magic
tech sky130A
magscale 1 2
timestamp 1763991652
<< obsli1 >>
rect 1104 2159 19228 20145
<< obsm1 >>
rect 934 2128 19288 20392
<< metal2 >>
rect 1582 21714 1638 22514
rect 2134 21714 2190 22514
rect 2686 21714 2742 22514
rect 3238 21714 3294 22514
rect 3790 21714 3846 22514
rect 4342 21714 4398 22514
rect 4894 21714 4950 22514
rect 5446 21714 5502 22514
rect 5998 21714 6054 22514
rect 6550 21714 6606 22514
rect 7102 21714 7158 22514
rect 7654 21714 7710 22514
rect 8206 21714 8262 22514
rect 8758 21714 8814 22514
rect 9310 21714 9366 22514
rect 9862 21714 9918 22514
rect 10414 21714 10470 22514
rect 10966 21714 11022 22514
rect 11518 21714 11574 22514
rect 12070 21714 12126 22514
rect 12622 21714 12678 22514
rect 13174 21714 13230 22514
rect 13726 21714 13782 22514
rect 14278 21714 14334 22514
rect 14830 21714 14886 22514
rect 15382 21714 15438 22514
rect 15934 21714 15990 22514
rect 16486 21714 16542 22514
rect 17038 21714 17094 22514
rect 17590 21714 17646 22514
rect 18142 21714 18198 22514
rect 18694 21714 18750 22514
rect 15198 0 15254 800
<< obsm2 >>
rect 938 21658 1526 21842
rect 1694 21658 2078 21842
rect 2246 21658 2630 21842
rect 2798 21658 3182 21842
rect 3350 21658 3734 21842
rect 3902 21658 4286 21842
rect 4454 21658 4838 21842
rect 5006 21658 5390 21842
rect 5558 21658 5942 21842
rect 6110 21658 6494 21842
rect 6662 21658 7046 21842
rect 7214 21658 7598 21842
rect 7766 21658 8150 21842
rect 8318 21658 8702 21842
rect 8870 21658 9254 21842
rect 9422 21658 9806 21842
rect 9974 21658 10358 21842
rect 10526 21658 10910 21842
rect 11078 21658 11462 21842
rect 11630 21658 12014 21842
rect 12182 21658 12566 21842
rect 12734 21658 13118 21842
rect 13286 21658 13670 21842
rect 13838 21658 14222 21842
rect 14390 21658 14774 21842
rect 14942 21658 15326 21842
rect 15494 21658 15878 21842
rect 16046 21658 16430 21842
rect 16598 21658 16982 21842
rect 17150 21658 17534 21842
rect 17702 21658 18086 21842
rect 18254 21658 18638 21842
rect 18806 21658 18932 21842
rect 938 856 18932 21658
rect 938 800 15142 856
rect 15310 800 18932 856
<< metal3 >>
rect 0 16600 800 16720
rect 19570 11160 20370 11280
rect 0 5448 800 5568
<< obsm3 >>
rect 800 16800 19570 20161
rect 880 16520 19570 16800
rect 800 11360 19570 16520
rect 800 11080 19490 11360
rect 800 5648 19570 11080
rect 880 5368 19570 5648
rect 800 2143 19570 5368
<< metal4 >>
rect 3209 2128 3529 20176
rect 3869 2128 4189 20176
rect 7740 2128 8060 20176
rect 8400 2128 8720 20176
rect 12271 2128 12591 20176
rect 12931 2128 13251 20176
rect 16802 2128 17122 20176
rect 17462 2128 17782 20176
<< obsm4 >>
rect 4291 8195 4357 12477
<< metal5 >>
rect 1056 18384 19276 18704
rect 1056 17724 19276 18044
rect 1056 13896 19276 14216
rect 1056 13236 19276 13556
rect 1056 9408 19276 9728
rect 1056 8748 19276 9068
rect 1056 4920 19276 5240
rect 1056 4260 19276 4580
<< labels >>
rlabel metal4 s 3869 2128 4189 20176 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8400 2128 8720 20176 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12931 2128 13251 20176 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17462 2128 17782 20176 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4920 19276 5240 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9408 19276 9728 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13896 19276 14216 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18384 19276 18704 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3209 2128 3529 20176 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7740 2128 8060 20176 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12271 2128 12591 20176 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16802 2128 17122 20176 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4260 19276 4580 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8748 19276 9068 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13236 19276 13556 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 17724 19276 18044 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 19570 11160 20370 11280 6 clk
port 3 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 p
port 4 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 rst
port 5 nsew signal input
rlabel metal2 s 1582 21714 1638 22514 6 x[0]
port 6 nsew signal input
rlabel metal2 s 7102 21714 7158 22514 6 x[10]
port 7 nsew signal input
rlabel metal2 s 7654 21714 7710 22514 6 x[11]
port 8 nsew signal input
rlabel metal2 s 8206 21714 8262 22514 6 x[12]
port 9 nsew signal input
rlabel metal2 s 8758 21714 8814 22514 6 x[13]
port 10 nsew signal input
rlabel metal2 s 9310 21714 9366 22514 6 x[14]
port 11 nsew signal input
rlabel metal2 s 9862 21714 9918 22514 6 x[15]
port 12 nsew signal input
rlabel metal2 s 10414 21714 10470 22514 6 x[16]
port 13 nsew signal input
rlabel metal2 s 10966 21714 11022 22514 6 x[17]
port 14 nsew signal input
rlabel metal2 s 11518 21714 11574 22514 6 x[18]
port 15 nsew signal input
rlabel metal2 s 12070 21714 12126 22514 6 x[19]
port 16 nsew signal input
rlabel metal2 s 2134 21714 2190 22514 6 x[1]
port 17 nsew signal input
rlabel metal2 s 12622 21714 12678 22514 6 x[20]
port 18 nsew signal input
rlabel metal2 s 13174 21714 13230 22514 6 x[21]
port 19 nsew signal input
rlabel metal2 s 13726 21714 13782 22514 6 x[22]
port 20 nsew signal input
rlabel metal2 s 14278 21714 14334 22514 6 x[23]
port 21 nsew signal input
rlabel metal2 s 14830 21714 14886 22514 6 x[24]
port 22 nsew signal input
rlabel metal2 s 15382 21714 15438 22514 6 x[25]
port 23 nsew signal input
rlabel metal2 s 15934 21714 15990 22514 6 x[26]
port 24 nsew signal input
rlabel metal2 s 16486 21714 16542 22514 6 x[27]
port 25 nsew signal input
rlabel metal2 s 17038 21714 17094 22514 6 x[28]
port 26 nsew signal input
rlabel metal2 s 17590 21714 17646 22514 6 x[29]
port 27 nsew signal input
rlabel metal2 s 2686 21714 2742 22514 6 x[2]
port 28 nsew signal input
rlabel metal2 s 18142 21714 18198 22514 6 x[30]
port 29 nsew signal input
rlabel metal2 s 18694 21714 18750 22514 6 x[31]
port 30 nsew signal input
rlabel metal2 s 3238 21714 3294 22514 6 x[3]
port 31 nsew signal input
rlabel metal2 s 3790 21714 3846 22514 6 x[4]
port 32 nsew signal input
rlabel metal2 s 4342 21714 4398 22514 6 x[5]
port 33 nsew signal input
rlabel metal2 s 4894 21714 4950 22514 6 x[6]
port 34 nsew signal input
rlabel metal2 s 5446 21714 5502 22514 6 x[7]
port 35 nsew signal input
rlabel metal2 s 5998 21714 6054 22514 6 x[8]
port 36 nsew signal input
rlabel metal2 s 6550 21714 6606 22514 6 x[9]
port 37 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 y
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20370 22514
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 977224
string GDS_FILE /openlane/designs/spm/runs/openlane_test/results/signoff/spm.magic.gds
string GDS_START 117684
<< end >>

