magic
tech sky130A
magscale 1 2
timestamp 1763991656
<< checkpaint >>
rect -1260 7244 21630 23774
rect -2866 -1260 21630 7244
<< viali >>
rect 5549 20009 5583 20043
rect 17325 20009 17359 20043
rect 3893 19941 3927 19975
rect 8493 19941 8527 19975
rect 15393 19941 15427 19975
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2789 19805 2823 19839
rect 3341 19805 3375 19839
rect 4077 19805 4111 19839
rect 4445 19805 4479 19839
rect 5181 19805 5215 19839
rect 5733 19805 5767 19839
rect 6561 19805 6595 19839
rect 6837 19805 6871 19839
rect 7389 19805 7423 19839
rect 7941 19805 7975 19839
rect 8309 19805 8343 19839
rect 9137 19805 9171 19839
rect 9597 19805 9631 19839
rect 9965 19805 9999 19839
rect 10517 19805 10551 19839
rect 11069 19805 11103 19839
rect 11621 19805 11655 19839
rect 12173 19805 12207 19839
rect 12725 19805 12759 19839
rect 13645 19805 13679 19839
rect 13921 19805 13955 19839
rect 14381 19805 14415 19839
rect 14565 19805 14599 19839
rect 14657 19805 14691 19839
rect 14933 19805 14967 19839
rect 15209 19805 15243 19839
rect 15485 19805 15519 19839
rect 16037 19805 16071 19839
rect 16865 19805 16899 19839
rect 16957 19805 16991 19839
rect 17049 19805 17083 19839
rect 17141 19805 17175 19839
rect 17509 19805 17543 19839
rect 17785 19805 17819 19839
rect 18061 19805 18095 19839
rect 18429 19805 18463 19839
rect 18889 19805 18923 19839
rect 1869 19669 1903 19703
rect 2421 19669 2455 19703
rect 2973 19669 3007 19703
rect 3525 19669 3559 19703
rect 4629 19669 4663 19703
rect 4997 19669 5031 19703
rect 6377 19669 6411 19703
rect 6653 19669 6687 19703
rect 7205 19669 7239 19703
rect 7757 19669 7791 19703
rect 8953 19669 8987 19703
rect 9413 19669 9447 19703
rect 10149 19669 10183 19703
rect 10701 19669 10735 19703
rect 11253 19669 11287 19703
rect 11805 19669 11839 19703
rect 12357 19669 12391 19703
rect 12909 19669 12943 19703
rect 13553 19669 13587 19703
rect 13737 19669 13771 19703
rect 14197 19669 14231 19703
rect 14841 19669 14875 19703
rect 15117 19669 15151 19703
rect 15669 19669 15703 19703
rect 16221 19669 16255 19703
rect 16681 19669 16715 19703
rect 17601 19669 17635 19703
rect 17877 19669 17911 19703
rect 18245 19669 18279 19703
rect 18705 19669 18739 19703
rect 8769 19465 8803 19499
rect 15025 19465 15059 19499
rect 10517 19397 10551 19431
rect 15577 19397 15611 19431
rect 16957 19397 16991 19431
rect 3617 19329 3651 19363
rect 4169 19329 4203 19363
rect 4445 19329 4479 19363
rect 7021 19329 7055 19363
rect 9229 19329 9263 19363
rect 9965 19329 9999 19363
rect 10425 19329 10459 19363
rect 10609 19329 10643 19363
rect 11713 19329 11747 19363
rect 12357 19329 12391 19363
rect 15209 19329 15243 19363
rect 15393 19329 15427 19363
rect 16681 19329 16715 19363
rect 2973 19261 3007 19295
rect 3065 19261 3099 19295
rect 3157 19261 3191 19295
rect 3249 19261 3283 19295
rect 4077 19261 4111 19295
rect 4721 19261 4755 19295
rect 7297 19261 7331 19295
rect 9321 19261 9355 19295
rect 10057 19261 10091 19295
rect 12633 19261 12667 19295
rect 14105 19261 14139 19295
rect 14381 19261 14415 19295
rect 16221 19261 16255 19295
rect 2789 19125 2823 19159
rect 3525 19125 3559 19159
rect 3893 19125 3927 19159
rect 6193 19125 6227 19159
rect 8861 19125 8895 19159
rect 10241 19125 10275 19159
rect 11621 19125 11655 19159
rect 15301 19125 15335 19159
rect 18429 19125 18463 19159
rect 4629 18921 4663 18955
rect 5181 18921 5215 18955
rect 8125 18921 8159 18955
rect 10590 18921 10624 18955
rect 13093 18921 13127 18955
rect 16681 18921 16715 18955
rect 17417 18921 17451 18955
rect 3617 18853 3651 18887
rect 14105 18853 14139 18887
rect 1869 18785 1903 18819
rect 3893 18785 3927 18819
rect 4537 18785 4571 18819
rect 4997 18785 5031 18819
rect 5365 18785 5399 18819
rect 5457 18785 5491 18819
rect 6653 18785 6687 18819
rect 7297 18785 7331 18819
rect 7757 18785 7791 18819
rect 8309 18785 8343 18819
rect 10057 18785 10091 18819
rect 10333 18785 10367 18819
rect 13277 18785 13311 18819
rect 13369 18785 13403 18819
rect 14381 18785 14415 18819
rect 14933 18785 14967 18819
rect 17601 18785 17635 18819
rect 17877 18785 17911 18819
rect 18337 18785 18371 18819
rect 1777 18717 1811 18751
rect 4813 18717 4847 18751
rect 5549 18717 5583 18751
rect 5641 18717 5675 18751
rect 5917 18717 5951 18751
rect 6561 18717 6595 18751
rect 7573 18717 7607 18751
rect 8401 18717 8435 18751
rect 8493 18717 8527 18751
rect 8585 18717 8619 18751
rect 8953 18717 8987 18751
rect 9597 18717 9631 18751
rect 9689 18717 9723 18751
rect 9873 18717 9907 18751
rect 13461 18717 13495 18751
rect 13553 18717 13587 18751
rect 14473 18717 14507 18751
rect 16957 18717 16991 18751
rect 17325 18717 17359 18751
rect 17969 18717 18003 18751
rect 2145 18649 2179 18683
rect 7389 18649 7423 18683
rect 15209 18649 15243 18683
rect 16865 18649 16899 18683
rect 1685 18581 1719 18615
rect 12081 18581 12115 18615
rect 18889 18581 18923 18615
rect 4721 18377 4755 18411
rect 5917 18377 5951 18411
rect 10701 18377 10735 18411
rect 15025 18377 15059 18411
rect 2881 18309 2915 18343
rect 3157 18241 3191 18275
rect 3617 18241 3651 18275
rect 4721 18241 4755 18275
rect 4905 18241 4939 18275
rect 6009 18241 6043 18275
rect 6745 18241 6779 18275
rect 8493 18241 8527 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9597 18241 9631 18275
rect 10333 18241 10367 18275
rect 11253 18241 11287 18275
rect 13277 18241 13311 18275
rect 13461 18241 13495 18275
rect 15393 18241 15427 18275
rect 18705 18241 18739 18275
rect 18889 18241 18923 18275
rect 3249 18173 3283 18207
rect 3525 18173 3559 18207
rect 6837 18173 6871 18207
rect 8585 18173 8619 18207
rect 9505 18173 9539 18207
rect 10241 18173 10275 18207
rect 10425 18173 10459 18207
rect 10517 18173 10551 18207
rect 15485 18173 15519 18207
rect 18521 18173 18555 18207
rect 6377 18105 6411 18139
rect 8861 18105 8895 18139
rect 1409 18037 1443 18071
rect 9045 18037 9079 18071
rect 10057 18037 10091 18071
rect 13369 18037 13403 18071
rect 7205 17833 7239 17867
rect 18521 17833 18555 17867
rect 10425 17697 10459 17731
rect 11897 17697 11931 17731
rect 12449 17697 12483 17731
rect 13277 17697 13311 17731
rect 16773 17697 16807 17731
rect 5457 17629 5491 17663
rect 10149 17629 10183 17663
rect 13369 17629 13403 17663
rect 15669 17629 15703 17663
rect 15853 17629 15887 17663
rect 5733 17561 5767 17595
rect 17049 17561 17083 17595
rect 13093 17493 13127 17527
rect 13737 17493 13771 17527
rect 15853 17493 15887 17527
rect 5917 17289 5951 17323
rect 11253 17289 11287 17323
rect 16313 17289 16347 17323
rect 17693 17289 17727 17323
rect 3249 17221 3283 17255
rect 13921 17221 13955 17255
rect 15577 17221 15611 17255
rect 1409 17153 1443 17187
rect 2329 17153 2363 17187
rect 2881 17153 2915 17187
rect 3157 17153 3191 17187
rect 3341 17153 3375 17187
rect 4813 17153 4847 17187
rect 4905 17153 4939 17187
rect 5535 17153 5569 17187
rect 5917 17159 5951 17193
rect 6101 17153 6135 17187
rect 8401 17153 8435 17187
rect 11161 17153 11195 17187
rect 12357 17153 12391 17187
rect 12817 17153 12851 17187
rect 12909 17153 12943 17187
rect 13645 17153 13679 17187
rect 15669 17153 15703 17187
rect 15945 17153 15979 17187
rect 17601 17153 17635 17187
rect 2973 17085 3007 17119
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 5365 17085 5399 17119
rect 8493 17085 8527 17119
rect 11989 17085 12023 17119
rect 12449 17085 12483 17119
rect 16037 17085 16071 17119
rect 5825 17017 5859 17051
rect 12633 17017 12667 17051
rect 1593 16949 1627 16983
rect 2237 16949 2271 16983
rect 2605 16949 2639 16983
rect 4629 16949 4663 16983
rect 8033 16949 8067 16983
rect 15393 16949 15427 16983
rect 6561 16745 6595 16779
rect 8953 16745 8987 16779
rect 10701 16745 10735 16779
rect 2881 16609 2915 16643
rect 4077 16609 4111 16643
rect 7573 16609 7607 16643
rect 7665 16609 7699 16643
rect 15761 16609 15795 16643
rect 15853 16609 15887 16643
rect 15945 16609 15979 16643
rect 16313 16609 16347 16643
rect 18061 16609 18095 16643
rect 18797 16609 18831 16643
rect 3157 16541 3191 16575
rect 3801 16541 3835 16575
rect 5641 16541 5675 16575
rect 6469 16541 6503 16575
rect 7757 16541 7791 16575
rect 7849 16541 7883 16575
rect 8125 16541 8159 16575
rect 8677 16541 8711 16575
rect 9505 16541 9539 16575
rect 16037 16541 16071 16575
rect 12173 16473 12207 16507
rect 16589 16473 16623 16507
rect 1409 16405 1443 16439
rect 5549 16405 5583 16439
rect 6285 16405 6319 16439
rect 7389 16405 7423 16439
rect 16221 16405 16255 16439
rect 18245 16405 18279 16439
rect 4537 16201 4571 16235
rect 8217 16201 8251 16235
rect 8309 16201 8343 16235
rect 8953 16201 8987 16235
rect 13277 16201 13311 16235
rect 17417 16201 17451 16235
rect 1869 16133 1903 16167
rect 5365 16133 5399 16167
rect 10425 16133 10459 16167
rect 17693 16133 17727 16167
rect 4629 16065 4663 16099
rect 5089 16065 5123 16099
rect 5549 16065 5583 16099
rect 5733 16065 5767 16099
rect 6469 16065 6503 16099
rect 8493 16065 8527 16099
rect 10701 16065 10735 16099
rect 10977 16065 11011 16099
rect 11529 16065 11563 16099
rect 13921 16065 13955 16099
rect 15669 16065 15703 16099
rect 17325 16065 17359 16099
rect 17877 16065 17911 16099
rect 18061 16065 18095 16099
rect 18521 16065 18555 16099
rect 5181 15997 5215 16031
rect 6745 15997 6779 16031
rect 8677 15997 8711 16031
rect 10885 15997 10919 16031
rect 11805 15997 11839 16031
rect 18613 15997 18647 16031
rect 11345 15929 11379 15963
rect 18153 15929 18187 15963
rect 2145 15861 2179 15895
rect 4721 15861 4755 15895
rect 13829 15861 13863 15895
rect 15577 15861 15611 15895
rect 7389 15657 7423 15691
rect 9873 15657 9907 15691
rect 11161 15657 11195 15691
rect 11989 15657 12023 15691
rect 8493 15589 8527 15623
rect 2237 15521 2271 15555
rect 2697 15521 2731 15555
rect 8033 15521 8067 15555
rect 8677 15521 8711 15555
rect 12173 15521 12207 15555
rect 13921 15521 13955 15555
rect 14565 15521 14599 15555
rect 15209 15521 15243 15555
rect 15669 15521 15703 15555
rect 2605 15453 2639 15487
rect 4353 15453 4387 15487
rect 7297 15453 7331 15487
rect 8125 15453 8159 15487
rect 8585 15453 8619 15487
rect 8769 15453 8803 15487
rect 9965 15453 9999 15487
rect 11069 15453 11103 15487
rect 11253 15453 11287 15487
rect 11897 15453 11931 15487
rect 15485 15453 15519 15487
rect 12449 15385 12483 15419
rect 3801 15317 3835 15351
rect 15301 15317 15335 15351
rect 3157 15113 3191 15147
rect 13093 15113 13127 15147
rect 7113 15045 7147 15079
rect 3433 14977 3467 15011
rect 3617 14977 3651 15011
rect 6745 14977 6779 15011
rect 7021 14977 7055 15011
rect 7205 14977 7239 15011
rect 10793 14977 10827 15011
rect 10885 14977 10919 15011
rect 13369 14977 13403 15011
rect 13737 14977 13771 15011
rect 13921 14977 13955 15011
rect 14473 14977 14507 15011
rect 15853 14977 15887 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 17509 14977 17543 15011
rect 1409 14909 1443 14943
rect 1685 14909 1719 14943
rect 6837 14909 6871 14943
rect 10701 14909 10735 14943
rect 10977 14909 11011 14943
rect 11529 14909 11563 14943
rect 12081 14909 12115 14943
rect 13277 14909 13311 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 14565 14909 14599 14943
rect 17601 14909 17635 14943
rect 3249 14841 3283 14875
rect 14105 14841 14139 14875
rect 6469 14773 6503 14807
rect 10517 14773 10551 14807
rect 13829 14773 13863 14807
rect 15945 14773 15979 14807
rect 16221 14773 16255 14807
rect 17141 14773 17175 14807
rect 2329 14569 2363 14603
rect 5549 14569 5583 14603
rect 7021 14569 7055 14603
rect 10136 14569 10170 14603
rect 12541 14569 12575 14603
rect 16773 14569 16807 14603
rect 18889 14569 18923 14603
rect 2145 14501 2179 14535
rect 2513 14433 2547 14467
rect 2789 14433 2823 14467
rect 4077 14433 4111 14467
rect 6561 14433 6595 14467
rect 7573 14433 7607 14467
rect 9873 14433 9907 14467
rect 11621 14433 11655 14467
rect 12357 14433 12391 14467
rect 12817 14433 12851 14467
rect 13461 14433 13495 14467
rect 15025 14433 15059 14467
rect 17141 14433 17175 14467
rect 2053 14365 2087 14399
rect 2605 14365 2639 14399
rect 2697 14365 2731 14399
rect 2973 14365 3007 14399
rect 3157 14365 3191 14399
rect 3801 14365 3835 14399
rect 5825 14365 5859 14399
rect 6653 14365 6687 14399
rect 6745 14365 6779 14399
rect 6837 14365 6871 14399
rect 9045 14365 9079 14399
rect 12909 14365 12943 14399
rect 13553 14365 13587 14399
rect 5733 14297 5767 14331
rect 15301 14297 15335 14331
rect 17417 14297 17451 14331
rect 3065 14229 3099 14263
rect 6377 14229 6411 14263
rect 9137 14229 9171 14263
rect 11805 14229 11839 14263
rect 13185 14229 13219 14263
rect 6101 14025 6135 14059
rect 10977 14025 11011 14059
rect 11529 14025 11563 14059
rect 15669 14025 15703 14059
rect 18521 14025 18555 14059
rect 4629 13957 4663 13991
rect 6653 13957 6687 13991
rect 14841 13957 14875 13991
rect 2421 13889 2455 13923
rect 6009 13889 6043 13923
rect 8309 13889 8343 13923
rect 10885 13889 10919 13923
rect 11713 13889 11747 13923
rect 11805 13889 11839 13923
rect 12909 13889 12943 13923
rect 14933 13889 14967 13923
rect 15853 13889 15887 13923
rect 16129 13889 16163 13923
rect 17969 13889 18003 13923
rect 18153 13889 18187 13923
rect 18429 13889 18463 13923
rect 2329 13821 2363 13855
rect 6377 13821 6411 13855
rect 13185 13821 13219 13855
rect 14657 13821 14691 13855
rect 15945 13821 15979 13855
rect 16037 13821 16071 13855
rect 17233 13821 17267 13855
rect 17877 13821 17911 13855
rect 18337 13821 18371 13855
rect 2697 13685 2731 13719
rect 4905 13685 4939 13719
rect 8125 13685 8159 13719
rect 8572 13685 8606 13719
rect 10057 13685 10091 13719
rect 6561 13481 6595 13515
rect 7113 13481 7147 13515
rect 12541 13481 12575 13515
rect 17141 13481 17175 13515
rect 4629 13345 4663 13379
rect 5089 13345 5123 13379
rect 7389 13345 7423 13379
rect 8677 13345 8711 13379
rect 10793 13345 10827 13379
rect 16957 13345 16991 13379
rect 3801 13277 3835 13311
rect 4997 13277 5031 13311
rect 7481 13277 7515 13311
rect 8953 13277 8987 13311
rect 9413 13277 9447 13311
rect 9597 13277 9631 13311
rect 9689 13277 9723 13311
rect 10241 13277 10275 13311
rect 16865 13277 16899 13311
rect 5273 13209 5307 13243
rect 11069 13209 11103 13243
rect 3893 13141 3927 13175
rect 8125 13141 8159 13175
rect 9045 13141 9079 13175
rect 9229 13141 9263 13175
rect 6193 12937 6227 12971
rect 7481 12937 7515 12971
rect 9689 12937 9723 12971
rect 11069 12937 11103 12971
rect 11805 12937 11839 12971
rect 14289 12937 14323 12971
rect 18889 12937 18923 12971
rect 4721 12869 4755 12903
rect 13001 12869 13035 12903
rect 2605 12801 2639 12835
rect 7665 12801 7699 12835
rect 7849 12801 7883 12835
rect 10149 12801 10183 12835
rect 10701 12801 10735 12835
rect 11713 12801 11747 12835
rect 15577 12801 15611 12835
rect 15945 12801 15979 12835
rect 16129 12801 16163 12835
rect 17141 12801 17175 12835
rect 4445 12733 4479 12767
rect 7941 12733 7975 12767
rect 8217 12733 8251 12767
rect 10057 12733 10091 12767
rect 10609 12733 10643 12767
rect 15485 12733 15519 12767
rect 15669 12733 15703 12767
rect 15761 12733 15795 12767
rect 17417 12733 17451 12767
rect 3893 12597 3927 12631
rect 9781 12597 9815 12631
rect 15301 12597 15335 12631
rect 16037 12597 16071 12631
rect 5641 12393 5675 12427
rect 7849 12393 7883 12427
rect 9781 12393 9815 12427
rect 11253 12393 11287 12427
rect 18429 12393 18463 12427
rect 17693 12325 17727 12359
rect 1409 12257 1443 12291
rect 3893 12257 3927 12291
rect 5733 12257 5767 12291
rect 14565 12257 14599 12291
rect 16037 12257 16071 12291
rect 16221 12257 16255 12291
rect 16957 12257 16991 12291
rect 17601 12257 17635 12291
rect 17969 12257 18003 12291
rect 6469 12189 6503 12223
rect 6837 12189 6871 12223
rect 8401 12189 8435 12223
rect 11161 12189 11195 12223
rect 11345 12189 11379 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 13829 12189 13863 12223
rect 14289 12189 14323 12223
rect 18061 12189 18095 12223
rect 18521 12189 18555 12223
rect 1685 12121 1719 12155
rect 4169 12121 4203 12155
rect 6561 12121 6595 12155
rect 11069 12121 11103 12155
rect 3157 12053 3191 12087
rect 6377 12053 6411 12087
rect 6929 12053 6963 12087
rect 12817 12053 12851 12087
rect 13277 12053 13311 12087
rect 16865 12053 16899 12087
rect 1961 11849 1995 11883
rect 2145 11849 2179 11883
rect 4261 11849 4295 11883
rect 8125 11849 8159 11883
rect 8953 11849 8987 11883
rect 13737 11849 13771 11883
rect 15393 11849 15427 11883
rect 15761 11849 15795 11883
rect 12265 11781 12299 11815
rect 1869 11713 1903 11747
rect 2329 11713 2363 11747
rect 2421 11713 2455 11747
rect 3893 11713 3927 11747
rect 4537 11713 4571 11747
rect 5825 11713 5859 11747
rect 6377 11713 6411 11747
rect 8401 11713 8435 11747
rect 9229 11713 9263 11747
rect 9321 11713 9355 11747
rect 9413 11713 9447 11747
rect 9597 11713 9631 11747
rect 9781 11713 9815 11747
rect 14197 11713 14231 11747
rect 15485 11713 15519 11747
rect 15945 11713 15979 11747
rect 16129 11713 16163 11747
rect 16865 11713 16899 11747
rect 2513 11645 2547 11679
rect 2605 11645 2639 11679
rect 2789 11645 2823 11679
rect 3341 11645 3375 11679
rect 3985 11645 4019 11679
rect 4445 11645 4479 11679
rect 4629 11645 4663 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 5549 11645 5583 11679
rect 5641 11645 5675 11679
rect 6009 11645 6043 11679
rect 6653 11645 6687 11679
rect 8309 11645 8343 11679
rect 9137 11645 9171 11679
rect 11989 11645 12023 11679
rect 14289 11645 14323 11679
rect 16773 11645 16807 11679
rect 17233 11645 17267 11679
rect 3525 11577 3559 11611
rect 8769 11577 8803 11611
rect 9689 11509 9723 11543
rect 13829 11509 13863 11543
rect 2605 11305 2639 11339
rect 6469 11305 6503 11339
rect 13461 11305 13495 11339
rect 12265 11237 12299 11271
rect 2973 11169 3007 11203
rect 6653 11169 6687 11203
rect 7113 11169 7147 11203
rect 10609 11169 10643 11203
rect 10701 11169 10735 11203
rect 12449 11169 12483 11203
rect 12633 11169 12667 11203
rect 2789 11101 2823 11135
rect 6745 11101 6779 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 10793 11101 10827 11135
rect 10885 11101 10919 11135
rect 12081 11101 12115 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 12909 11101 12943 11135
rect 13093 11101 13127 11135
rect 13553 11101 13587 11135
rect 18337 11101 18371 11135
rect 10425 10965 10459 10999
rect 11529 10965 11563 10999
rect 13001 10965 13035 10999
rect 18889 10965 18923 10999
rect 4445 10761 4479 10795
rect 11069 10761 11103 10795
rect 11529 10761 11563 10795
rect 18429 10761 18463 10795
rect 9597 10693 9631 10727
rect 11253 10693 11287 10727
rect 15577 10693 15611 10727
rect 3985 10625 4019 10659
rect 4997 10625 5031 10659
rect 5181 10625 5215 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 7757 10625 7791 10659
rect 11337 10625 11371 10659
rect 11713 10625 11747 10659
rect 12541 10625 12575 10659
rect 15209 10625 15243 10659
rect 15485 10625 15519 10659
rect 15669 10625 15703 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 4077 10557 4111 10591
rect 7941 10557 7975 10591
rect 9321 10557 9355 10591
rect 11897 10557 11931 10591
rect 12449 10557 12483 10591
rect 15301 10557 15335 10591
rect 16681 10557 16715 10591
rect 16957 10557 16991 10591
rect 12909 10489 12943 10523
rect 4261 10421 4295 10455
rect 5273 10421 5307 10455
rect 7573 10421 7607 10455
rect 14933 10421 14967 10455
rect 18521 10421 18555 10455
rect 3985 10217 4019 10251
rect 5917 10217 5951 10251
rect 10517 10217 10551 10251
rect 11989 10217 12023 10251
rect 12541 10217 12575 10251
rect 16589 10217 16623 10251
rect 17693 10217 17727 10251
rect 16129 10149 16163 10183
rect 3157 10081 3191 10115
rect 4169 10081 4203 10115
rect 4445 10081 4479 10115
rect 6653 10081 6687 10115
rect 6745 10081 6779 10115
rect 7665 10081 7699 10115
rect 10977 10081 11011 10115
rect 14381 10081 14415 10115
rect 14657 10081 14691 10115
rect 16773 10081 16807 10115
rect 17877 10081 17911 10115
rect 18153 10081 18187 10115
rect 3249 10013 3283 10047
rect 3433 10013 3467 10047
rect 3893 10013 3927 10047
rect 4077 10013 4111 10047
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 7113 10013 7147 10047
rect 8401 10013 8435 10047
rect 8953 10013 8987 10047
rect 10885 10013 10919 10047
rect 11437 10013 11471 10047
rect 13277 10013 13311 10047
rect 16405 10013 16439 10047
rect 16865 10013 16899 10047
rect 16957 10013 16991 10047
rect 17049 10013 17083 10047
rect 17601 10013 17635 10047
rect 18245 10013 18279 10047
rect 2881 9945 2915 9979
rect 12265 9945 12299 9979
rect 16313 9945 16347 9979
rect 1409 9877 1443 9911
rect 3249 9877 3283 9911
rect 6469 9877 6503 9911
rect 7849 9877 7883 9911
rect 9045 9877 9079 9911
rect 13829 9877 13863 9911
rect 2145 9673 2179 9707
rect 2881 9673 2915 9707
rect 11529 9673 11563 9707
rect 18429 9673 18463 9707
rect 5917 9605 5951 9639
rect 9413 9605 9447 9639
rect 18613 9605 18647 9639
rect 2053 9527 2087 9561
rect 2513 9537 2547 9571
rect 4905 9537 4939 9571
rect 6193 9537 6227 9571
rect 6929 9537 6963 9571
rect 7205 9537 7239 9571
rect 7757 9537 7791 9571
rect 11161 9537 11195 9571
rect 11345 9537 11379 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 14657 9537 14691 9571
rect 14749 9537 14783 9571
rect 15025 9537 15059 9571
rect 16681 9537 16715 9571
rect 18521 9537 18555 9571
rect 2421 9469 2455 9503
rect 6561 9469 6595 9503
rect 7021 9469 7055 9503
rect 9689 9469 9723 9503
rect 12173 9469 12207 9503
rect 12449 9469 12483 9503
rect 12725 9469 12759 9503
rect 14381 9469 14415 9503
rect 16957 9469 16991 9503
rect 7941 9401 7975 9435
rect 5089 9333 5123 9367
rect 11253 9333 11287 9367
rect 12265 9333 12299 9367
rect 12909 9333 12943 9367
rect 8033 9129 8067 9163
rect 12633 9129 12667 9163
rect 13369 9129 13403 9163
rect 14657 9129 14691 9163
rect 16129 9129 16163 9163
rect 1961 8993 1995 9027
rect 2421 8993 2455 9027
rect 6285 8993 6319 9027
rect 11161 8993 11195 9027
rect 13645 8993 13679 9027
rect 14473 8993 14507 9027
rect 15945 8993 15979 9027
rect 2053 8925 2087 8959
rect 2513 8925 2547 8959
rect 9045 8925 9079 8959
rect 9321 8925 9355 8959
rect 11069 8925 11103 8959
rect 13277 8925 13311 8959
rect 13737 8925 13771 8959
rect 14289 8925 14323 8959
rect 14749 8925 14783 8959
rect 15853 8925 15887 8959
rect 6561 8857 6595 8891
rect 14105 8857 14139 8891
rect 3157 8789 3191 8823
rect 10701 8789 10735 8823
rect 7021 8585 7055 8619
rect 10885 8585 10919 8619
rect 13277 8585 13311 8619
rect 14657 8585 14691 8619
rect 4077 8517 4111 8551
rect 9413 8517 9447 8551
rect 11805 8517 11839 8551
rect 2697 8449 2731 8483
rect 3525 8449 3559 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4261 8449 4295 8483
rect 6929 8449 6963 8483
rect 9137 8449 9171 8483
rect 13369 8449 13403 8483
rect 15209 8449 15243 8483
rect 16037 8449 16071 8483
rect 16221 8449 16255 8483
rect 16681 8449 16715 8483
rect 2329 8381 2363 8415
rect 2789 8381 2823 8415
rect 2881 8381 2915 8415
rect 2973 8381 3007 8415
rect 3433 8381 3467 8415
rect 4537 8381 4571 8415
rect 11529 8381 11563 8415
rect 15485 8381 15519 8415
rect 16129 8381 16163 8415
rect 16313 8381 16347 8415
rect 16497 8381 16531 8415
rect 16957 8381 16991 8415
rect 2513 8313 2547 8347
rect 3893 8313 3927 8347
rect 1777 8245 1811 8279
rect 6009 8245 6043 8279
rect 18429 8245 18463 8279
rect 1777 8041 1811 8075
rect 4445 8041 4479 8075
rect 9505 8041 9539 8075
rect 10885 8041 10919 8075
rect 15853 8041 15887 8075
rect 17417 8041 17451 8075
rect 17601 8041 17635 8075
rect 7849 7973 7883 8007
rect 12357 7973 12391 8007
rect 1409 7905 1443 7939
rect 4813 7905 4847 7939
rect 8125 7905 8159 7939
rect 13553 7905 13587 7939
rect 14749 7905 14783 7939
rect 15025 7905 15059 7939
rect 18061 7905 18095 7939
rect 18337 7905 18371 7939
rect 1593 7837 1627 7871
rect 3617 7837 3651 7871
rect 4353 7837 4387 7871
rect 4905 7837 4939 7871
rect 4997 7837 5031 7871
rect 5089 7837 5123 7871
rect 7113 7837 7147 7871
rect 8217 7837 8251 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 9413 7837 9447 7871
rect 10333 7837 10367 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 15117 7837 15151 7871
rect 15209 7837 15243 7871
rect 15301 7837 15335 7871
rect 15485 7837 15519 7871
rect 15669 7837 15703 7871
rect 15761 7837 15795 7871
rect 15945 7837 15979 7871
rect 17325 7837 17359 7871
rect 17969 7837 18003 7871
rect 5273 7769 5307 7803
rect 7021 7769 7055 7803
rect 8585 7769 8619 7803
rect 13921 7769 13955 7803
rect 2329 7701 2363 7735
rect 4629 7701 4663 7735
rect 7757 7701 7791 7735
rect 9689 7701 9723 7735
rect 14841 7701 14875 7735
rect 15485 7701 15519 7735
rect 18889 7701 18923 7735
rect 1409 7497 1443 7531
rect 7021 7497 7055 7531
rect 10149 7497 10183 7531
rect 13645 7497 13679 7531
rect 18521 7497 18555 7531
rect 2881 7429 2915 7463
rect 4445 7429 4479 7463
rect 10333 7429 10367 7463
rect 3157 7361 3191 7395
rect 4169 7361 4203 7395
rect 6745 7361 6779 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 7941 7361 7975 7395
rect 9965 7361 9999 7395
rect 10241 7361 10275 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 11897 7361 11931 7395
rect 14933 7361 14967 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 18705 7361 18739 7395
rect 18889 7361 18923 7395
rect 5917 7293 5951 7327
rect 6653 7293 6687 7327
rect 8217 7293 8251 7327
rect 9781 7293 9815 7327
rect 12173 7293 12207 7327
rect 14105 7293 14139 7327
rect 14657 7293 14691 7327
rect 14841 7293 14875 7327
rect 15301 7293 15335 7327
rect 9689 7225 9723 7259
rect 6377 7157 6411 7191
rect 10425 7157 10459 7191
rect 16773 7157 16807 7191
rect 2329 6953 2363 6987
rect 4169 6953 4203 6987
rect 9045 6953 9079 6987
rect 12909 6953 12943 6987
rect 14197 6953 14231 6987
rect 9321 6817 9355 6851
rect 15393 6817 15427 6851
rect 16129 6817 16163 6851
rect 17877 6817 17911 6851
rect 2237 6749 2271 6783
rect 2973 6749 3007 6783
rect 3157 6749 3191 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 8953 6749 8987 6783
rect 9505 6749 9539 6783
rect 11621 6749 11655 6783
rect 12081 6749 12115 6783
rect 12265 6749 12299 6783
rect 12817 6749 12851 6783
rect 14749 6749 14783 6783
rect 15301 6749 15335 6783
rect 15577 6749 15611 6783
rect 16037 6749 16071 6783
rect 16221 6749 16255 6783
rect 16313 6749 16347 6783
rect 16589 6749 16623 6783
rect 17141 6749 17175 6783
rect 3893 6681 3927 6715
rect 11989 6681 12023 6715
rect 3157 6613 3191 6647
rect 9689 6613 9723 6647
rect 12265 6613 12299 6647
rect 14933 6613 14967 6647
rect 15669 6613 15703 6647
rect 15853 6613 15887 6647
rect 17325 6613 17359 6647
rect 18889 6409 18923 6443
rect 7389 6341 7423 6375
rect 16681 6341 16715 6375
rect 17417 6341 17451 6375
rect 3157 6273 3191 6307
rect 3617 6273 3651 6307
rect 4537 6273 4571 6307
rect 4721 6273 4755 6307
rect 7113 6273 7147 6307
rect 9873 6273 9907 6307
rect 10609 6273 10643 6307
rect 11897 6273 11931 6307
rect 14565 6273 14599 6307
rect 16865 6273 16899 6307
rect 16957 6273 16991 6307
rect 17141 6273 17175 6307
rect 2881 6205 2915 6239
rect 3709 6205 3743 6239
rect 8861 6205 8895 6239
rect 8953 6205 8987 6239
rect 11713 6205 11747 6239
rect 11805 6205 11839 6239
rect 11989 6205 12023 6239
rect 12173 6205 12207 6239
rect 12817 6205 12851 6239
rect 14841 6205 14875 6239
rect 3249 6137 3283 6171
rect 16313 6137 16347 6171
rect 1409 6069 1443 6103
rect 4629 6069 4663 6103
rect 9597 6069 9631 6103
rect 9689 6069 9723 6103
rect 10701 6069 10735 6103
rect 11529 6069 11563 6103
rect 2329 5865 2363 5899
rect 8217 5865 8251 5899
rect 9505 5865 9539 5899
rect 9952 5865 9986 5899
rect 13001 5865 13035 5899
rect 17049 5865 17083 5899
rect 18337 5865 18371 5899
rect 7389 5797 7423 5831
rect 11437 5797 11471 5831
rect 15853 5797 15887 5831
rect 2789 5729 2823 5763
rect 2881 5729 2915 5763
rect 4445 5729 4479 5763
rect 5365 5729 5399 5763
rect 5549 5729 5583 5763
rect 5917 5729 5951 5763
rect 8493 5729 8527 5763
rect 9321 5729 9355 5763
rect 9689 5729 9723 5763
rect 12449 5729 12483 5763
rect 13369 5729 13403 5763
rect 16313 5729 16347 5763
rect 16681 5729 16715 5763
rect 1501 5661 1535 5695
rect 2237 5661 2271 5695
rect 2697 5661 2731 5695
rect 2973 5661 3007 5695
rect 4537 5661 4571 5695
rect 5089 5661 5123 5695
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 5641 5661 5675 5695
rect 8125 5661 8159 5695
rect 8585 5661 8619 5695
rect 9137 5661 9171 5695
rect 9413 5661 9447 5695
rect 11621 5661 11655 5695
rect 12541 5661 12575 5695
rect 13185 5661 13219 5695
rect 16228 5661 16262 5695
rect 16773 5661 16807 5695
rect 18429 5661 18463 5695
rect 8953 5593 8987 5627
rect 1593 5525 1627 5559
rect 2513 5525 2547 5559
rect 4905 5525 4939 5559
rect 7481 5525 7515 5559
rect 12265 5525 12299 5559
rect 12909 5525 12943 5559
rect 3157 5321 3191 5355
rect 6745 5321 6779 5355
rect 10701 5321 10735 5355
rect 14013 5321 14047 5355
rect 15945 5321 15979 5355
rect 4721 5253 4755 5287
rect 9229 5253 9263 5287
rect 12541 5253 12575 5287
rect 3341 5185 3375 5219
rect 6653 5185 6687 5219
rect 8401 5185 8435 5219
rect 8953 5185 8987 5219
rect 11897 5185 11931 5219
rect 12265 5185 12299 5219
rect 14197 5185 14231 5219
rect 3525 5117 3559 5151
rect 3617 5117 3651 5151
rect 4169 5117 4203 5151
rect 4445 5117 4479 5151
rect 8585 5117 8619 5151
rect 11529 5117 11563 5151
rect 11989 5117 12023 5151
rect 14473 5117 14507 5151
rect 6193 4981 6227 5015
rect 3801 4777 3835 4811
rect 5733 4777 5767 4811
rect 9505 4777 9539 4811
rect 13369 4777 13403 4811
rect 15117 4777 15151 4811
rect 3525 4709 3559 4743
rect 1777 4641 1811 4675
rect 2053 4641 2087 4675
rect 4261 4641 4295 4675
rect 4169 4573 4203 4607
rect 5825 4573 5859 4607
rect 9413 4573 9447 4607
rect 13277 4573 13311 4607
rect 15025 4573 15059 4607
rect 2789 4233 2823 4267
rect 15025 4233 15059 4267
rect 15301 4165 15335 4199
rect 2697 4097 2731 4131
rect 15485 2601 15519 2635
rect 15301 2397 15335 2431
<< metal1 >>
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 17494 20380 17500 20392
rect 16632 20352 17500 20380
rect 16632 20340 16638 20352
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 1104 20154 19228 20176
rect 1104 20102 3215 20154
rect 3267 20102 3279 20154
rect 3331 20102 3343 20154
rect 3395 20102 3407 20154
rect 3459 20102 3471 20154
rect 3523 20102 7746 20154
rect 7798 20102 7810 20154
rect 7862 20102 7874 20154
rect 7926 20102 7938 20154
rect 7990 20102 8002 20154
rect 8054 20102 12277 20154
rect 12329 20102 12341 20154
rect 12393 20102 12405 20154
rect 12457 20102 12469 20154
rect 12521 20102 12533 20154
rect 12585 20102 16808 20154
rect 16860 20102 16872 20154
rect 16924 20102 16936 20154
rect 16988 20102 17000 20154
rect 17052 20102 17064 20154
rect 17116 20102 19228 20154
rect 1104 20080 19228 20102
rect 3142 20000 3148 20052
rect 3200 20040 3206 20052
rect 5537 20043 5595 20049
rect 5537 20040 5549 20043
rect 3200 20012 5549 20040
rect 3200 20000 3206 20012
rect 5537 20009 5549 20012
rect 5583 20009 5595 20043
rect 5537 20003 5595 20009
rect 6546 20000 6552 20052
rect 6604 20000 6610 20052
rect 13814 20000 13820 20052
rect 13872 20000 13878 20052
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 17862 20040 17868 20052
rect 17359 20012 17868 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 2958 19932 2964 19984
rect 3016 19972 3022 19984
rect 3881 19975 3939 19981
rect 3881 19972 3893 19975
rect 3016 19944 3893 19972
rect 3016 19932 3022 19944
rect 3881 19941 3893 19944
rect 3927 19941 3939 19975
rect 3881 19935 3939 19941
rect 6564 19904 6592 20000
rect 8481 19975 8539 19981
rect 8481 19941 8493 19975
rect 8527 19972 8539 19975
rect 9214 19972 9220 19984
rect 8527 19944 9220 19972
rect 8527 19941 8539 19944
rect 8481 19935 8539 19941
rect 9214 19932 9220 19944
rect 9272 19932 9278 19984
rect 13832 19972 13860 20000
rect 15381 19975 15439 19981
rect 13832 19944 14688 19972
rect 6564 19876 6868 19904
rect 1578 19796 1584 19848
rect 1636 19836 1642 19848
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1636 19808 1685 19836
rect 1636 19796 1642 19808
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 2130 19796 2136 19848
rect 2188 19836 2194 19848
rect 2225 19839 2283 19845
rect 2225 19836 2237 19839
rect 2188 19808 2237 19836
rect 2188 19796 2194 19808
rect 2225 19805 2237 19808
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2774 19796 2780 19848
rect 2832 19796 2838 19848
rect 3050 19796 3056 19848
rect 3108 19836 3114 19848
rect 3329 19839 3387 19845
rect 3329 19836 3341 19839
rect 3108 19808 3341 19836
rect 3108 19796 3114 19808
rect 3329 19805 3341 19808
rect 3375 19805 3387 19839
rect 3329 19799 3387 19805
rect 3786 19796 3792 19848
rect 3844 19836 3850 19848
rect 4065 19839 4123 19845
rect 4065 19836 4077 19839
rect 3844 19808 4077 19836
rect 3844 19796 3850 19808
rect 4065 19805 4077 19808
rect 4111 19805 4123 19839
rect 4065 19799 4123 19805
rect 4338 19796 4344 19848
rect 4396 19836 4402 19848
rect 4433 19839 4491 19845
rect 4433 19836 4445 19839
rect 4396 19808 4445 19836
rect 4396 19796 4402 19808
rect 4433 19805 4445 19808
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 4948 19808 5181 19836
rect 4948 19796 4954 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 5534 19796 5540 19848
rect 5592 19836 5598 19848
rect 5721 19839 5779 19845
rect 5721 19836 5733 19839
rect 5592 19808 5733 19836
rect 5592 19796 5598 19808
rect 5721 19805 5733 19808
rect 5767 19805 5779 19839
rect 5721 19799 5779 19805
rect 5994 19796 6000 19848
rect 6052 19836 6058 19848
rect 6840 19845 6868 19876
rect 13170 19864 13176 19916
rect 13228 19904 13234 19916
rect 13228 19876 13952 19904
rect 13228 19864 13234 19876
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 6052 19808 6561 19836
rect 6052 19796 6058 19808
rect 6549 19805 6561 19808
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 7156 19808 7389 19836
rect 7156 19796 7162 19808
rect 7377 19805 7389 19808
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 7650 19796 7656 19848
rect 7708 19836 7714 19848
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 7708 19808 7941 19836
rect 7708 19796 7714 19808
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 8294 19796 8300 19848
rect 8352 19796 8358 19848
rect 8754 19796 8760 19848
rect 8812 19836 8818 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 8812 19808 9137 19836
rect 8812 19796 8818 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 9585 19839 9643 19845
rect 9585 19836 9597 19839
rect 9364 19808 9597 19836
rect 9364 19796 9370 19808
rect 9585 19805 9597 19808
rect 9631 19805 9643 19839
rect 9585 19799 9643 19805
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9916 19808 9965 19836
rect 9916 19796 9922 19808
rect 9953 19805 9965 19808
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 10410 19796 10416 19848
rect 10468 19836 10474 19848
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 10468 19808 10517 19836
rect 10468 19796 10474 19808
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 11054 19796 11060 19848
rect 11112 19796 11118 19848
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 11609 19839 11667 19845
rect 11609 19836 11621 19839
rect 11572 19808 11621 19836
rect 11572 19796 11578 19808
rect 11609 19805 11621 19808
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 12124 19808 12173 19836
rect 12124 19796 12130 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 13924 19845 13952 19876
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12676 19808 12725 19836
rect 12676 19796 12682 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19805 13967 19839
rect 13909 19799 13967 19805
rect 13648 19768 13676 19799
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 14366 19796 14372 19848
rect 14424 19796 14430 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 14660 19845 14688 19944
rect 15381 19941 15393 19975
rect 15427 19972 15439 19975
rect 15746 19972 15752 19984
rect 15427 19944 15752 19972
rect 15427 19941 15439 19944
rect 15381 19935 15439 19941
rect 15746 19932 15752 19944
rect 15804 19932 15810 19984
rect 17954 19972 17960 19984
rect 17144 19944 17960 19972
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 14292 19768 14320 19796
rect 14936 19768 14964 19799
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 15436 19808 15485 19836
rect 15436 19796 15442 19808
rect 15473 19805 15485 19808
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15988 19808 16037 19836
rect 15988 19796 15994 19808
rect 16025 19805 16037 19808
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 17144 19845 17172 19944
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 17218 19864 17224 19916
rect 17276 19864 17282 19916
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 17644 19876 18092 19904
rect 17644 19864 17650 19876
rect 16853 19839 16911 19845
rect 16853 19836 16865 19839
rect 16632 19808 16865 19836
rect 16632 19796 16638 19808
rect 16853 19805 16865 19808
rect 16899 19805 16911 19839
rect 16853 19799 16911 19805
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 16960 19768 16988 19799
rect 2976 19740 3648 19768
rect 13648 19740 14044 19768
rect 14292 19740 14964 19768
rect 15028 19740 16988 19768
rect 1854 19660 1860 19712
rect 1912 19660 1918 19712
rect 2130 19660 2136 19712
rect 2188 19700 2194 19712
rect 2976 19709 3004 19740
rect 2409 19703 2467 19709
rect 2409 19700 2421 19703
rect 2188 19672 2421 19700
rect 2188 19660 2194 19672
rect 2409 19669 2421 19672
rect 2455 19669 2467 19703
rect 2409 19663 2467 19669
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19669 3019 19703
rect 2961 19663 3019 19669
rect 3510 19660 3516 19712
rect 3568 19660 3574 19712
rect 3620 19700 3648 19740
rect 14016 19712 14044 19740
rect 4522 19700 4528 19712
rect 3620 19672 4528 19700
rect 4522 19660 4528 19672
rect 4580 19660 4586 19712
rect 4614 19660 4620 19712
rect 4672 19660 4678 19712
rect 4982 19660 4988 19712
rect 5040 19660 5046 19712
rect 6362 19660 6368 19712
rect 6420 19660 6426 19712
rect 6546 19660 6552 19712
rect 6604 19700 6610 19712
rect 6641 19703 6699 19709
rect 6641 19700 6653 19703
rect 6604 19672 6653 19700
rect 6604 19660 6610 19672
rect 6641 19669 6653 19672
rect 6687 19669 6699 19703
rect 6641 19663 6699 19669
rect 7190 19660 7196 19712
rect 7248 19660 7254 19712
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7432 19672 7757 19700
rect 7432 19660 7438 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 8938 19660 8944 19712
rect 8996 19660 9002 19712
rect 9398 19660 9404 19712
rect 9456 19660 9462 19712
rect 10134 19660 10140 19712
rect 10192 19660 10198 19712
rect 10689 19703 10747 19709
rect 10689 19669 10701 19703
rect 10735 19700 10747 19703
rect 10778 19700 10784 19712
rect 10735 19672 10784 19700
rect 10735 19669 10747 19672
rect 10689 19663 10747 19669
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 11238 19660 11244 19712
rect 11296 19660 11302 19712
rect 11790 19660 11796 19712
rect 11848 19660 11854 19712
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 11940 19672 12357 19700
rect 11940 19660 11946 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 12345 19663 12403 19669
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19700 12955 19703
rect 13446 19700 13452 19712
rect 12943 19672 13452 19700
rect 12943 19669 12955 19672
rect 12897 19663 12955 19669
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 13630 19700 13636 19712
rect 13587 19672 13636 19700
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 13722 19660 13728 19712
rect 13780 19660 13786 19712
rect 13998 19660 14004 19712
rect 14056 19660 14062 19712
rect 14182 19660 14188 19712
rect 14240 19660 14246 19712
rect 14829 19703 14887 19709
rect 14829 19669 14841 19703
rect 14875 19700 14887 19703
rect 15028 19700 15056 19740
rect 15396 19712 15424 19740
rect 14875 19672 15056 19700
rect 14875 19669 14887 19672
rect 14829 19663 14887 19669
rect 15102 19660 15108 19712
rect 15160 19660 15166 19712
rect 15378 19660 15384 19712
rect 15436 19660 15442 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15528 19672 15669 19700
rect 15528 19660 15534 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15657 19663 15715 19669
rect 16206 19660 16212 19712
rect 16264 19660 16270 19712
rect 16666 19660 16672 19712
rect 16724 19660 16730 19712
rect 17052 19700 17080 19799
rect 17236 19768 17264 19864
rect 17494 19796 17500 19848
rect 17552 19796 17558 19848
rect 18064 19845 18092 19876
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 17788 19768 17816 19799
rect 18138 19796 18144 19848
rect 18196 19836 18202 19848
rect 18417 19839 18475 19845
rect 18417 19836 18429 19839
rect 18196 19808 18429 19836
rect 18196 19796 18202 19808
rect 18417 19805 18429 19808
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18748 19808 18889 19836
rect 18748 19796 18754 19808
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 17236 19740 17816 19768
rect 17310 19700 17316 19712
rect 17052 19672 17316 19700
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 17589 19703 17647 19709
rect 17589 19700 17601 19703
rect 17460 19672 17601 19700
rect 17460 19660 17466 19672
rect 17589 19669 17601 19672
rect 17635 19669 17647 19703
rect 17589 19663 17647 19669
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 17865 19703 17923 19709
rect 17865 19700 17877 19703
rect 17736 19672 17877 19700
rect 17736 19660 17742 19672
rect 17865 19669 17877 19672
rect 17911 19669 17923 19703
rect 17865 19663 17923 19669
rect 18230 19660 18236 19712
rect 18288 19660 18294 19712
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 1104 19610 19228 19632
rect 1104 19558 3875 19610
rect 3927 19558 3939 19610
rect 3991 19558 4003 19610
rect 4055 19558 4067 19610
rect 4119 19558 4131 19610
rect 4183 19558 8406 19610
rect 8458 19558 8470 19610
rect 8522 19558 8534 19610
rect 8586 19558 8598 19610
rect 8650 19558 8662 19610
rect 8714 19558 12937 19610
rect 12989 19558 13001 19610
rect 13053 19558 13065 19610
rect 13117 19558 13129 19610
rect 13181 19558 13193 19610
rect 13245 19558 17468 19610
rect 17520 19558 17532 19610
rect 17584 19558 17596 19610
rect 17648 19558 17660 19610
rect 17712 19558 17724 19610
rect 17776 19558 19228 19610
rect 1104 19536 19228 19558
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 8803 19468 9260 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 9030 19428 9036 19440
rect 8510 19400 9036 19428
rect 9030 19388 9036 19400
rect 9088 19388 9094 19440
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 2832 19332 3617 19360
rect 2832 19320 2838 19332
rect 3605 19329 3617 19332
rect 3651 19360 3663 19363
rect 3878 19360 3884 19372
rect 3651 19332 3884 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 3878 19320 3884 19332
rect 3936 19320 3942 19372
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2924 19264 2973 19292
rect 2924 19252 2930 19264
rect 2961 19261 2973 19264
rect 3007 19261 3019 19295
rect 2961 19255 3019 19261
rect 3050 19252 3056 19304
rect 3108 19252 3114 19304
rect 3145 19295 3203 19301
rect 3145 19261 3157 19295
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 3970 19292 3976 19304
rect 3283 19264 3976 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 2590 19184 2596 19236
rect 2648 19224 2654 19236
rect 3160 19224 3188 19255
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19261 4123 19295
rect 4172 19292 4200 19323
rect 4246 19320 4252 19372
rect 4304 19360 4310 19372
rect 4433 19363 4491 19369
rect 4433 19360 4445 19363
rect 4304 19332 4445 19360
rect 4304 19320 4310 19332
rect 4433 19329 4445 19332
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 5810 19320 5816 19372
rect 5868 19320 5874 19372
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 9232 19369 9260 19468
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10318 19496 10324 19508
rect 10192 19468 10324 19496
rect 10192 19456 10198 19468
rect 10318 19456 10324 19468
rect 10376 19496 10382 19508
rect 10376 19468 10640 19496
rect 10376 19456 10382 19468
rect 10505 19431 10563 19437
rect 10505 19428 10517 19431
rect 9968 19400 10517 19428
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6880 19332 7021 19360
rect 6880 19320 6886 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9766 19360 9772 19372
rect 9263 19332 9772 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 9968 19369 9996 19400
rect 10505 19397 10517 19400
rect 10551 19397 10563 19431
rect 10505 19391 10563 19397
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10612 19369 10640 19468
rect 14366 19456 14372 19508
rect 14424 19456 14430 19508
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 15013 19499 15071 19505
rect 15013 19496 15025 19499
rect 14608 19468 15025 19496
rect 14608 19456 14614 19468
rect 15013 19465 15025 19468
rect 15059 19465 15071 19499
rect 15013 19459 15071 19465
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 16724 19468 16988 19496
rect 16724 19456 16730 19468
rect 11054 19388 11060 19440
rect 11112 19428 11118 19440
rect 11112 19400 12388 19428
rect 11112 19388 11118 19400
rect 10413 19363 10471 19369
rect 10413 19360 10425 19363
rect 10192 19332 10425 19360
rect 10192 19320 10198 19332
rect 10413 19329 10425 19332
rect 10459 19329 10471 19363
rect 10413 19323 10471 19329
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 11330 19320 11336 19372
rect 11388 19360 11394 19372
rect 12360 19369 12388 19400
rect 13630 19388 13636 19440
rect 13688 19388 13694 19440
rect 14384 19428 14412 19456
rect 16960 19437 16988 19468
rect 15565 19431 15623 19437
rect 15565 19428 15577 19431
rect 14384 19400 15577 19428
rect 15565 19397 15577 19400
rect 15611 19397 15623 19431
rect 15565 19391 15623 19397
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19397 17003 19431
rect 16945 19391 17003 19397
rect 17402 19388 17408 19440
rect 17460 19388 17466 19440
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11388 19332 11713 19360
rect 11388 19320 11394 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 4338 19292 4344 19304
rect 4172 19264 4344 19292
rect 4065 19255 4123 19261
rect 4080 19224 4108 19255
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4706 19252 4712 19304
rect 4764 19252 4770 19304
rect 7282 19252 7288 19304
rect 7340 19252 7346 19304
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19292 9367 19295
rect 9674 19292 9680 19304
rect 9355 19264 9680 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 10045 19295 10103 19301
rect 10045 19261 10057 19295
rect 10091 19292 10103 19295
rect 11146 19292 11152 19304
rect 10091 19264 11152 19292
rect 10091 19261 10103 19264
rect 10045 19255 10103 19261
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 12618 19252 12624 19304
rect 12676 19252 12682 19304
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14139 19264 14381 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14369 19261 14381 19264
rect 14415 19261 14427 19295
rect 15212 19292 15240 19323
rect 15378 19320 15384 19372
rect 15436 19320 15442 19372
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 16209 19295 16267 19301
rect 15212 19264 15424 19292
rect 14369 19255 14427 19261
rect 4430 19224 4436 19236
rect 2648 19196 2912 19224
rect 3160 19196 4016 19224
rect 4080 19196 4436 19224
rect 2648 19184 2654 19196
rect 2774 19116 2780 19168
rect 2832 19116 2838 19168
rect 2884 19156 2912 19196
rect 3513 19159 3571 19165
rect 3513 19156 3525 19159
rect 2884 19128 3525 19156
rect 3513 19125 3525 19128
rect 3559 19125 3571 19159
rect 3513 19119 3571 19125
rect 3786 19116 3792 19168
rect 3844 19156 3850 19168
rect 3881 19159 3939 19165
rect 3881 19156 3893 19159
rect 3844 19128 3893 19156
rect 3844 19116 3850 19128
rect 3881 19125 3893 19128
rect 3927 19125 3939 19159
rect 3988 19156 4016 19196
rect 4430 19184 4436 19196
rect 4488 19184 4494 19236
rect 15396 19168 15424 19264
rect 16209 19261 16221 19295
rect 16255 19292 16267 19295
rect 16255 19264 16344 19292
rect 16255 19261 16267 19264
rect 16209 19255 16267 19261
rect 16316 19168 16344 19264
rect 4890 19156 4896 19168
rect 3988 19128 4896 19156
rect 3881 19119 3939 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 6178 19116 6184 19168
rect 6236 19116 6242 19168
rect 8846 19116 8852 19168
rect 8904 19116 8910 19168
rect 10226 19116 10232 19168
rect 10284 19116 10290 19168
rect 11606 19116 11612 19168
rect 11664 19116 11670 19168
rect 15286 19116 15292 19168
rect 15344 19116 15350 19168
rect 15378 19116 15384 19168
rect 15436 19116 15442 19168
rect 16298 19116 16304 19168
rect 16356 19116 16362 19168
rect 18414 19116 18420 19168
rect 18472 19116 18478 19168
rect 1104 19066 19228 19088
rect 1104 19014 3215 19066
rect 3267 19014 3279 19066
rect 3331 19014 3343 19066
rect 3395 19014 3407 19066
rect 3459 19014 3471 19066
rect 3523 19014 7746 19066
rect 7798 19014 7810 19066
rect 7862 19014 7874 19066
rect 7926 19014 7938 19066
rect 7990 19014 8002 19066
rect 8054 19014 12277 19066
rect 12329 19014 12341 19066
rect 12393 19014 12405 19066
rect 12457 19014 12469 19066
rect 12521 19014 12533 19066
rect 12585 19014 16808 19066
rect 16860 19014 16872 19066
rect 16924 19014 16936 19066
rect 16988 19014 17000 19066
rect 17052 19014 17064 19066
rect 17116 19014 19228 19066
rect 1104 18992 19228 19014
rect 2682 18952 2688 18964
rect 1780 18924 2688 18952
rect 1780 18757 1808 18924
rect 2682 18912 2688 18924
rect 2740 18912 2746 18964
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 4617 18955 4675 18961
rect 4617 18952 4629 18955
rect 4028 18924 4629 18952
rect 4028 18912 4034 18924
rect 4617 18921 4629 18924
rect 4663 18921 4675 18955
rect 4617 18915 4675 18921
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 5169 18955 5227 18961
rect 5169 18952 5181 18955
rect 4764 18924 5181 18952
rect 4764 18912 4770 18924
rect 5169 18921 5181 18924
rect 5215 18921 5227 18955
rect 5169 18915 5227 18921
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7340 18924 8125 18952
rect 7340 18912 7346 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 8846 18912 8852 18964
rect 8904 18912 8910 18964
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 10134 18952 10140 18964
rect 9364 18924 10140 18952
rect 9364 18912 9370 18924
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 10578 18955 10636 18961
rect 10578 18952 10590 18955
rect 10284 18924 10590 18952
rect 10284 18912 10290 18924
rect 10578 18921 10590 18924
rect 10624 18921 10636 18955
rect 10578 18915 10636 18921
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 13081 18955 13139 18961
rect 13081 18952 13093 18955
rect 12676 18924 13093 18952
rect 12676 18912 12682 18924
rect 13081 18921 13093 18924
rect 13127 18921 13139 18955
rect 16298 18952 16304 18964
rect 13081 18915 13139 18921
rect 14384 18924 16304 18952
rect 3605 18887 3663 18893
rect 3605 18853 3617 18887
rect 3651 18884 3663 18887
rect 3694 18884 3700 18896
rect 3651 18856 3700 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 3694 18844 3700 18856
rect 3752 18884 3758 18896
rect 3752 18856 3924 18884
rect 3752 18844 3758 18856
rect 3896 18825 3924 18856
rect 4430 18844 4436 18896
rect 4488 18884 4494 18896
rect 5534 18884 5540 18896
rect 4488 18856 5396 18884
rect 4488 18844 4494 18856
rect 5368 18828 5396 18856
rect 5460 18856 5540 18884
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 3881 18819 3939 18825
rect 1903 18788 3188 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 3160 18760 3188 18788
rect 3881 18785 3893 18819
rect 3927 18785 3939 18819
rect 3881 18779 3939 18785
rect 4525 18819 4583 18825
rect 4525 18785 4537 18819
rect 4571 18816 4583 18819
rect 4985 18819 5043 18825
rect 4985 18816 4997 18819
rect 4571 18788 4997 18816
rect 4571 18785 4583 18788
rect 4525 18779 4583 18785
rect 4985 18785 4997 18788
rect 5031 18785 5043 18819
rect 4985 18779 5043 18785
rect 5350 18776 5356 18828
rect 5408 18776 5414 18828
rect 5460 18825 5488 18856
rect 5534 18844 5540 18856
rect 5592 18884 5598 18896
rect 6362 18884 6368 18896
rect 5592 18856 6368 18884
rect 5592 18844 5598 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 5445 18819 5503 18825
rect 5445 18785 5457 18819
rect 5491 18785 5503 18819
rect 5445 18779 5503 18785
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 6638 18816 6644 18828
rect 6236 18788 6644 18816
rect 6236 18776 6242 18788
rect 6638 18776 6644 18788
rect 6696 18776 6702 18828
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7331 18788 7757 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 8297 18819 8355 18825
rect 8297 18785 8309 18819
rect 8343 18816 8355 18819
rect 8864 18816 8892 18912
rect 14093 18887 14151 18893
rect 14093 18884 14105 18887
rect 13280 18856 14105 18884
rect 13280 18828 13308 18856
rect 14093 18853 14105 18856
rect 14139 18853 14151 18887
rect 14093 18847 14151 18853
rect 8343 18788 8892 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 9824 18788 10057 18816
rect 9824 18776 9830 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 10134 18776 10140 18828
rect 10192 18816 10198 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 10192 18788 10333 18816
rect 10192 18776 10198 18788
rect 10321 18785 10333 18788
rect 10367 18816 10379 18819
rect 10962 18816 10968 18828
rect 10367 18788 10968 18816
rect 10367 18785 10379 18788
rect 10321 18779 10379 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 13262 18776 13268 18828
rect 13320 18776 13326 18828
rect 13357 18819 13415 18825
rect 13357 18785 13369 18819
rect 13403 18816 13415 18819
rect 13722 18816 13728 18828
rect 13403 18788 13728 18816
rect 13403 18785 13415 18788
rect 13357 18779 13415 18785
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 14182 18776 14188 18828
rect 14240 18776 14246 18828
rect 14384 18825 14412 18924
rect 16298 18912 16304 18924
rect 16356 18952 16362 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16356 18924 16681 18952
rect 16356 18912 16362 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 16669 18915 16727 18921
rect 17402 18912 17408 18964
rect 17460 18912 17466 18964
rect 16574 18844 16580 18896
rect 16632 18884 16638 18896
rect 18506 18884 18512 18896
rect 16632 18856 16804 18884
rect 16632 18844 16638 18856
rect 16776 18828 16804 18856
rect 17880 18856 18512 18884
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18816 14979 18819
rect 14967 18788 16712 18816
rect 14967 18785 14979 18788
rect 14921 18779 14979 18785
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 3142 18708 3148 18760
rect 3200 18708 3206 18760
rect 4430 18708 4436 18760
rect 4488 18748 4494 18760
rect 4801 18751 4859 18757
rect 4801 18748 4813 18751
rect 4488 18720 4813 18748
rect 4488 18708 4494 18720
rect 4801 18717 4813 18720
rect 4847 18717 4859 18751
rect 4801 18711 4859 18717
rect 4890 18708 4896 18760
rect 4948 18748 4954 18760
rect 5537 18751 5595 18757
rect 5537 18748 5549 18751
rect 4948 18720 5549 18748
rect 4948 18708 4954 18720
rect 5537 18717 5549 18720
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18748 5687 18751
rect 5905 18751 5963 18757
rect 5905 18748 5917 18751
rect 5675 18720 5917 18748
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 5905 18717 5917 18720
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 6549 18751 6607 18757
rect 6549 18717 6561 18751
rect 6595 18717 6607 18751
rect 6549 18711 6607 18717
rect 2133 18683 2191 18689
rect 2133 18649 2145 18683
rect 2179 18649 2191 18683
rect 2133 18643 2191 18649
rect 1673 18615 1731 18621
rect 1673 18581 1685 18615
rect 1719 18612 1731 18615
rect 1762 18612 1768 18624
rect 1719 18584 1768 18612
rect 1719 18581 1731 18584
rect 1673 18575 1731 18581
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 2148 18612 2176 18643
rect 2590 18640 2596 18692
rect 2648 18640 2654 18692
rect 3878 18640 3884 18692
rect 3936 18680 3942 18692
rect 5994 18680 6000 18692
rect 3936 18652 6000 18680
rect 3936 18640 3942 18652
rect 5994 18640 6000 18652
rect 6052 18640 6058 18692
rect 6564 18680 6592 18711
rect 7558 18708 7564 18760
rect 7616 18708 7622 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 7377 18683 7435 18689
rect 7377 18680 7389 18683
rect 6564 18652 7389 18680
rect 7377 18649 7389 18652
rect 7423 18649 7435 18683
rect 8404 18680 8432 18711
rect 8478 18708 8484 18760
rect 8536 18708 8542 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8619 18720 8953 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18748 9643 18751
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 9631 18720 9689 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 9677 18717 9689 18720
rect 9723 18717 9735 18751
rect 9677 18711 9735 18717
rect 9858 18708 9864 18760
rect 9916 18708 9922 18760
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 13449 18751 13507 18757
rect 11664 18720 11730 18748
rect 11664 18708 11670 18720
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 14200 18748 14228 18776
rect 13587 18720 14228 18748
rect 14461 18751 14519 18757
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 14550 18748 14556 18760
rect 14507 18720 14556 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 9398 18680 9404 18692
rect 8404 18652 9404 18680
rect 7377 18643 7435 18649
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 13464 18680 13492 18711
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 13464 18652 13584 18680
rect 13556 18624 13584 18652
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 14936 18680 14964 18779
rect 16684 18760 16712 18788
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17880 18825 17908 18856
rect 18506 18844 18512 18856
rect 18564 18844 18570 18896
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 16816 18788 17601 18816
rect 16816 18776 16822 18788
rect 17589 18785 17601 18788
rect 17635 18785 17647 18819
rect 17589 18779 17647 18785
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18785 17923 18819
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 17865 18779 17923 18785
rect 17972 18788 18337 18816
rect 16666 18708 16672 18760
rect 16724 18708 16730 18760
rect 17972 18757 18000 18788
rect 18325 18785 18337 18788
rect 18371 18816 18383 18819
rect 18414 18816 18420 18828
rect 18371 18788 18420 18816
rect 18371 18785 18383 18788
rect 18325 18779 18383 18785
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18748 17003 18751
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 16991 18720 17325 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 13688 18652 14964 18680
rect 13688 18640 13694 18652
rect 15194 18640 15200 18692
rect 15252 18640 15258 18692
rect 16853 18683 16911 18689
rect 16853 18680 16865 18683
rect 16422 18652 16865 18680
rect 16853 18649 16865 18652
rect 16899 18649 16911 18683
rect 16853 18643 16911 18649
rect 2774 18612 2780 18624
rect 2148 18584 2780 18612
rect 2774 18572 2780 18584
rect 2832 18572 2838 18624
rect 8478 18572 8484 18624
rect 8536 18612 8542 18624
rect 10410 18612 10416 18624
rect 8536 18584 10416 18612
rect 8536 18572 8542 18584
rect 10410 18572 10416 18584
rect 10468 18572 10474 18624
rect 12066 18572 12072 18624
rect 12124 18572 12130 18624
rect 13538 18572 13544 18624
rect 13596 18572 13602 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 16960 18612 16988 18711
rect 16632 18584 16988 18612
rect 18877 18615 18935 18621
rect 16632 18572 16638 18584
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 18923 18584 19288 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 1104 18522 19228 18544
rect 1104 18470 3875 18522
rect 3927 18470 3939 18522
rect 3991 18470 4003 18522
rect 4055 18470 4067 18522
rect 4119 18470 4131 18522
rect 4183 18470 8406 18522
rect 8458 18470 8470 18522
rect 8522 18470 8534 18522
rect 8586 18470 8598 18522
rect 8650 18470 8662 18522
rect 8714 18470 12937 18522
rect 12989 18470 13001 18522
rect 13053 18470 13065 18522
rect 13117 18470 13129 18522
rect 13181 18470 13193 18522
rect 13245 18470 17468 18522
rect 17520 18470 17532 18522
rect 17584 18470 17596 18522
rect 17648 18470 17660 18522
rect 17712 18470 17724 18522
rect 17776 18470 19228 18522
rect 1104 18448 19228 18470
rect 3786 18408 3792 18420
rect 2884 18380 3792 18408
rect 2884 18349 2912 18380
rect 3786 18368 3792 18380
rect 3844 18368 3850 18420
rect 4338 18368 4344 18420
rect 4396 18408 4402 18420
rect 4709 18411 4767 18417
rect 4709 18408 4721 18411
rect 4396 18380 4721 18408
rect 4396 18368 4402 18380
rect 4709 18377 4721 18380
rect 4755 18377 4767 18411
rect 4709 18371 4767 18377
rect 5534 18368 5540 18420
rect 5592 18368 5598 18420
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 5905 18411 5963 18417
rect 5905 18408 5917 18411
rect 5868 18380 5917 18408
rect 5868 18368 5874 18380
rect 5905 18377 5917 18380
rect 5951 18377 5963 18411
rect 5905 18371 5963 18377
rect 6638 18368 6644 18420
rect 6696 18368 6702 18420
rect 9398 18368 9404 18420
rect 9456 18368 9462 18420
rect 9674 18368 9680 18420
rect 9732 18368 9738 18420
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 9916 18380 10701 18408
rect 9916 18368 9922 18380
rect 10689 18377 10701 18380
rect 10735 18377 10747 18411
rect 10689 18371 10747 18377
rect 13722 18368 13728 18420
rect 13780 18368 13786 18420
rect 15013 18411 15071 18417
rect 15013 18377 15025 18411
rect 15059 18408 15071 18411
rect 15194 18408 15200 18420
rect 15059 18380 15200 18408
rect 15059 18377 15071 18380
rect 15013 18371 15071 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 2869 18343 2927 18349
rect 2869 18309 2881 18343
rect 2915 18309 2927 18343
rect 4246 18340 4252 18352
rect 2869 18303 2927 18309
rect 3344 18312 4252 18340
rect 1762 18232 1768 18284
rect 1820 18232 1826 18284
rect 3142 18232 3148 18284
rect 3200 18272 3206 18284
rect 3344 18272 3372 18312
rect 3804 18284 3832 18312
rect 4246 18300 4252 18312
rect 4304 18300 4310 18352
rect 3200 18244 3372 18272
rect 3605 18275 3663 18281
rect 3200 18232 3206 18244
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 3694 18272 3700 18284
rect 3651 18244 3700 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 3786 18232 3792 18284
rect 3844 18232 3850 18284
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 4893 18275 4951 18281
rect 4755 18244 4844 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 2866 18164 2872 18216
rect 2924 18204 2930 18216
rect 3237 18207 3295 18213
rect 3237 18204 3249 18207
rect 2924 18176 3249 18204
rect 2924 18164 2930 18176
rect 3237 18173 3249 18176
rect 3283 18173 3295 18207
rect 3513 18207 3571 18213
rect 3513 18204 3525 18207
rect 3237 18167 3295 18173
rect 3344 18176 3525 18204
rect 1397 18071 1455 18077
rect 1397 18037 1409 18071
rect 1443 18068 1455 18071
rect 3344 18068 3372 18176
rect 3513 18173 3525 18176
rect 3559 18204 3571 18207
rect 4430 18204 4436 18216
rect 3559 18176 4436 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 4430 18164 4436 18176
rect 4488 18164 4494 18216
rect 4816 18080 4844 18244
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 5552 18272 5580 18368
rect 4939 18244 5580 18272
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 5994 18232 6000 18284
rect 6052 18232 6058 18284
rect 6656 18272 6684 18368
rect 9306 18340 9312 18352
rect 6932 18312 9312 18340
rect 6932 18284 6960 18312
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6656 18244 6745 18272
rect 6733 18241 6745 18244
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 6914 18232 6920 18284
rect 6972 18232 6978 18284
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 5350 18164 5356 18216
rect 5408 18164 5414 18216
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7558 18204 7564 18216
rect 6871 18176 7564 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 5368 18136 5396 18164
rect 6365 18139 6423 18145
rect 6365 18136 6377 18139
rect 5368 18108 6377 18136
rect 6365 18105 6377 18108
rect 6411 18105 6423 18139
rect 6365 18099 6423 18105
rect 1443 18040 3372 18068
rect 1443 18037 1455 18040
rect 1397 18031 1455 18037
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 5902 18068 5908 18080
rect 4856 18040 5908 18068
rect 4856 18028 4862 18040
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 8496 18068 8524 18235
rect 8846 18232 8852 18284
rect 8904 18232 8910 18284
rect 8956 18281 8984 18312
rect 9306 18300 9312 18312
rect 9364 18300 9370 18352
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18272 9183 18275
rect 9416 18272 9444 18368
rect 9692 18340 9720 18368
rect 12066 18340 12072 18352
rect 9692 18312 12072 18340
rect 9171 18244 9444 18272
rect 9585 18275 9643 18281
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9950 18272 9956 18284
rect 9631 18244 9956 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9950 18232 9956 18244
rect 10008 18272 10014 18284
rect 10008 18244 10180 18272
rect 10008 18232 10014 18244
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 8864 18204 8892 18232
rect 8619 18176 8892 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 9088 18176 9505 18204
rect 9088 18164 9094 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18136 8907 18139
rect 9674 18136 9680 18148
rect 8895 18108 9680 18136
rect 8895 18105 8907 18108
rect 8849 18099 8907 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8496 18040 9045 18068
rect 9033 18037 9045 18040
rect 9079 18037 9091 18071
rect 9033 18031 9091 18037
rect 10042 18028 10048 18080
rect 10100 18028 10106 18080
rect 10152 18068 10180 18244
rect 10318 18232 10324 18284
rect 10376 18232 10382 18284
rect 11256 18281 11284 18312
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18241 11299 18275
rect 11241 18235 11299 18241
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18272 13507 18275
rect 13740 18272 13768 18368
rect 13495 18244 13768 18272
rect 15304 18272 15332 18368
rect 18506 18300 18512 18352
rect 18564 18340 18570 18352
rect 18564 18312 18736 18340
rect 18564 18300 18570 18312
rect 18708 18281 18736 18312
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 15304 18244 15393 18272
rect 13495 18241 13507 18244
rect 13449 18235 13507 18241
rect 15381 18241 15393 18244
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18241 18751 18275
rect 18693 18235 18751 18241
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18272 18935 18275
rect 19260 18272 19288 18584
rect 18923 18244 19288 18272
rect 18923 18241 18935 18244
rect 18877 18235 18935 18241
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 10244 18136 10272 18167
rect 10410 18164 10416 18216
rect 10468 18164 10474 18216
rect 10505 18207 10563 18213
rect 10505 18173 10517 18207
rect 10551 18204 10563 18207
rect 11054 18204 11060 18216
rect 10551 18176 11060 18204
rect 10551 18173 10563 18176
rect 10505 18167 10563 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11974 18164 11980 18216
rect 12032 18164 12038 18216
rect 11146 18136 11152 18148
rect 10244 18108 11152 18136
rect 11146 18096 11152 18108
rect 11204 18136 11210 18148
rect 11992 18136 12020 18164
rect 11204 18108 12020 18136
rect 13280 18136 13308 18235
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18204 15531 18207
rect 16758 18204 16764 18216
rect 15519 18176 16764 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18012 18176 18521 18204
rect 18012 18164 18018 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 15378 18136 15384 18148
rect 13280 18108 15384 18136
rect 11204 18096 11210 18108
rect 15378 18096 15384 18108
rect 15436 18136 15442 18148
rect 15436 18108 15884 18136
rect 15436 18096 15442 18108
rect 15856 18080 15884 18108
rect 11330 18068 11336 18080
rect 10152 18040 11336 18068
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 13354 18028 13360 18080
rect 13412 18028 13418 18080
rect 15838 18028 15844 18080
rect 15896 18028 15902 18080
rect 1104 17978 19228 18000
rect 1104 17926 3215 17978
rect 3267 17926 3279 17978
rect 3331 17926 3343 17978
rect 3395 17926 3407 17978
rect 3459 17926 3471 17978
rect 3523 17926 7746 17978
rect 7798 17926 7810 17978
rect 7862 17926 7874 17978
rect 7926 17926 7938 17978
rect 7990 17926 8002 17978
rect 8054 17926 12277 17978
rect 12329 17926 12341 17978
rect 12393 17926 12405 17978
rect 12457 17926 12469 17978
rect 12521 17926 12533 17978
rect 12585 17926 16808 17978
rect 16860 17926 16872 17978
rect 16924 17926 16936 17978
rect 16988 17926 17000 17978
rect 17052 17926 17064 17978
rect 17116 17926 19228 17978
rect 1104 17904 19228 17926
rect 7193 17867 7251 17873
rect 7193 17833 7205 17867
rect 7239 17864 7251 17867
rect 7558 17864 7564 17876
rect 7239 17836 7564 17864
rect 7239 17833 7251 17836
rect 7193 17827 7251 17833
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 10042 17824 10048 17876
rect 10100 17824 10106 17876
rect 18506 17824 18512 17876
rect 18564 17824 18570 17876
rect 10060 17728 10088 17824
rect 10413 17731 10471 17737
rect 10413 17728 10425 17731
rect 10060 17700 10425 17728
rect 10413 17697 10425 17700
rect 10459 17697 10471 17731
rect 10413 17691 10471 17697
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12342 17728 12348 17740
rect 11931 17700 12348 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 12342 17688 12348 17700
rect 12400 17728 12406 17740
rect 12437 17731 12495 17737
rect 12437 17728 12449 17731
rect 12400 17700 12449 17728
rect 12400 17688 12406 17700
rect 12437 17697 12449 17700
rect 12483 17697 12495 17731
rect 12437 17691 12495 17697
rect 13262 17688 13268 17740
rect 13320 17688 13326 17740
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 16761 17731 16819 17737
rect 16761 17728 16773 17731
rect 16724 17700 16773 17728
rect 16724 17688 16730 17700
rect 16761 17697 16773 17700
rect 16807 17697 16819 17731
rect 16761 17691 16819 17697
rect 2866 17620 2872 17672
rect 2924 17660 2930 17672
rect 3050 17660 3056 17672
rect 2924 17632 3056 17660
rect 2924 17620 2930 17632
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3786 17620 3792 17672
rect 3844 17660 3850 17672
rect 5445 17663 5503 17669
rect 5445 17660 5457 17663
rect 3844 17632 5457 17660
rect 3844 17620 3850 17632
rect 5445 17629 5457 17632
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 10134 17620 10140 17672
rect 10192 17620 10198 17672
rect 13354 17620 13360 17672
rect 13412 17620 13418 17672
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15160 17632 15669 17660
rect 15160 17620 15166 17632
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 15896 17632 16160 17660
rect 15896 17620 15902 17632
rect 5718 17552 5724 17604
rect 5776 17552 5782 17604
rect 6454 17552 6460 17604
rect 6512 17552 6518 17604
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 16132 17536 16160 17632
rect 17034 17552 17040 17604
rect 17092 17552 17098 17604
rect 18046 17552 18052 17604
rect 18104 17552 18110 17604
rect 12802 17484 12808 17536
rect 12860 17524 12866 17536
rect 13081 17527 13139 17533
rect 13081 17524 13093 17527
rect 12860 17496 13093 17524
rect 12860 17484 12866 17496
rect 13081 17493 13093 17496
rect 13127 17493 13139 17527
rect 13081 17487 13139 17493
rect 13722 17484 13728 17536
rect 13780 17484 13786 17536
rect 15838 17484 15844 17536
rect 15896 17484 15902 17536
rect 16114 17484 16120 17536
rect 16172 17484 16178 17536
rect 1104 17434 19228 17456
rect 1104 17382 3875 17434
rect 3927 17382 3939 17434
rect 3991 17382 4003 17434
rect 4055 17382 4067 17434
rect 4119 17382 4131 17434
rect 4183 17382 8406 17434
rect 8458 17382 8470 17434
rect 8522 17382 8534 17434
rect 8586 17382 8598 17434
rect 8650 17382 8662 17434
rect 8714 17382 12937 17434
rect 12989 17382 13001 17434
rect 13053 17382 13065 17434
rect 13117 17382 13129 17434
rect 13181 17382 13193 17434
rect 13245 17382 17468 17434
rect 17520 17382 17532 17434
rect 17584 17382 17596 17434
rect 17648 17382 17660 17434
rect 17712 17382 17724 17434
rect 17776 17382 19228 17434
rect 1104 17360 19228 17382
rect 2682 17280 2688 17332
rect 2740 17280 2746 17332
rect 3142 17280 3148 17332
rect 3200 17320 3206 17332
rect 4798 17320 4804 17332
rect 3200 17292 3372 17320
rect 3200 17280 3206 17292
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 992 17156 1409 17184
rect 992 17144 998 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 2038 17144 2044 17196
rect 2096 17184 2102 17196
rect 2317 17187 2375 17193
rect 2317 17184 2329 17187
rect 2096 17156 2329 17184
rect 2096 17144 2102 17156
rect 2317 17153 2329 17156
rect 2363 17184 2375 17187
rect 2700 17184 2728 17280
rect 3237 17255 3295 17261
rect 3237 17252 3249 17255
rect 2884 17224 3249 17252
rect 2884 17193 2912 17224
rect 3237 17221 3249 17224
rect 3283 17221 3295 17255
rect 3237 17215 3295 17221
rect 3344 17193 3372 17292
rect 4632 17292 4804 17320
rect 2363 17156 2728 17184
rect 2869 17187 2927 17193
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 4632 17184 4660 17292
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 5905 17323 5963 17329
rect 5905 17320 5917 17323
rect 5828 17292 5917 17320
rect 5074 17252 5080 17264
rect 4816 17224 5080 17252
rect 4816 17193 4844 17224
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 3329 17147 3387 17153
rect 3436 17156 4660 17184
rect 4801 17187 4859 17193
rect 2682 17076 2688 17128
rect 2740 17076 2746 17128
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3050 17116 3056 17128
rect 3007 17088 3056 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 3160 17116 3188 17147
rect 3436 17116 3464 17156
rect 4801 17153 4813 17187
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17184 4951 17187
rect 5523 17187 5581 17193
rect 4939 17156 5488 17184
rect 4939 17153 4951 17156
rect 4893 17147 4951 17153
rect 3160 17088 3464 17116
rect 4985 17119 5043 17125
rect 4985 17085 4997 17119
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17116 5135 17119
rect 5258 17116 5264 17128
rect 5123 17088 5264 17116
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 2700 17048 2728 17076
rect 2700 17020 4844 17048
rect 1578 16940 1584 16992
rect 1636 16940 1642 16992
rect 2222 16940 2228 16992
rect 2280 16940 2286 16992
rect 2593 16983 2651 16989
rect 2593 16949 2605 16983
rect 2639 16980 2651 16983
rect 2866 16980 2872 16992
rect 2639 16952 2872 16980
rect 2639 16949 2651 16952
rect 2593 16943 2651 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 4614 16940 4620 16992
rect 4672 16940 4678 16992
rect 4816 16980 4844 17020
rect 4890 16980 4896 16992
rect 4816 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16980 4954 16992
rect 5000 16980 5028 17079
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5460 17116 5488 17156
rect 5523 17153 5535 17187
rect 5569 17184 5581 17187
rect 5828 17184 5856 17292
rect 5905 17289 5917 17292
rect 5951 17289 5963 17323
rect 5905 17283 5963 17289
rect 6546 17280 6552 17332
rect 6604 17280 6610 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11241 17323 11299 17329
rect 11241 17320 11253 17323
rect 11204 17292 11253 17320
rect 11204 17280 11210 17292
rect 11241 17289 11253 17292
rect 11287 17289 11299 17323
rect 11241 17283 11299 17289
rect 12342 17280 12348 17332
rect 12400 17280 12406 17332
rect 12802 17280 12808 17332
rect 12860 17280 12866 17332
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 13780 17292 13952 17320
rect 13780 17280 13786 17292
rect 5905 17196 5963 17199
rect 5569 17156 5856 17184
rect 5569 17153 5581 17156
rect 5523 17147 5581 17153
rect 5902 17144 5908 17196
rect 5960 17190 5966 17196
rect 5960 17162 5999 17190
rect 6089 17187 6147 17193
rect 5960 17144 5966 17162
rect 6089 17153 6101 17187
rect 6135 17184 6147 17187
rect 6564 17184 6592 17280
rect 11330 17212 11336 17264
rect 11388 17212 11394 17264
rect 6135 17156 6592 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 5460 17088 5948 17116
rect 5353 17079 5411 17085
rect 5368 17048 5396 17079
rect 5092 17020 5396 17048
rect 5092 16992 5120 17020
rect 5718 17008 5724 17060
rect 5776 17048 5782 17060
rect 5813 17051 5871 17057
rect 5813 17048 5825 17051
rect 5776 17020 5825 17048
rect 5776 17008 5782 17020
rect 5813 17017 5825 17020
rect 5859 17017 5871 17051
rect 5920 17048 5948 17088
rect 6196 17048 6224 17156
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8389 17187 8447 17193
rect 8389 17184 8401 17187
rect 8352 17156 8401 17184
rect 8352 17144 8358 17156
rect 8389 17153 8401 17156
rect 8435 17153 8447 17187
rect 8389 17147 8447 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11348 17184 11376 17212
rect 12360 17193 12388 17280
rect 12820 17252 12848 17280
rect 13924 17261 13952 17292
rect 15838 17280 15844 17332
rect 15896 17280 15902 17332
rect 16301 17323 16359 17329
rect 16301 17289 16313 17323
rect 16347 17320 16359 17323
rect 17034 17320 17040 17332
rect 16347 17292 17040 17320
rect 16347 17289 16359 17292
rect 16301 17283 16359 17289
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 17681 17323 17739 17329
rect 17681 17289 17693 17323
rect 17727 17320 17739 17323
rect 18046 17320 18052 17332
rect 17727 17292 18052 17320
rect 17727 17289 17739 17292
rect 17681 17283 17739 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 13909 17255 13967 17261
rect 12820 17224 12940 17252
rect 11195 17156 11376 17184
rect 12345 17187 12403 17193
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 12345 17153 12357 17187
rect 12391 17153 12403 17187
rect 12802 17184 12808 17196
rect 12345 17147 12403 17153
rect 12452 17156 12808 17184
rect 8478 17076 8484 17128
rect 8536 17076 8542 17128
rect 11974 17076 11980 17128
rect 12032 17076 12038 17128
rect 12452 17125 12480 17156
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 12912 17193 12940 17224
rect 13909 17221 13921 17255
rect 13955 17221 13967 17255
rect 15565 17255 15623 17261
rect 15565 17252 15577 17255
rect 15134 17224 15577 17252
rect 13909 17215 13967 17221
rect 15565 17221 15577 17224
rect 15611 17221 15623 17255
rect 15565 17215 15623 17221
rect 12897 17187 12955 17193
rect 12897 17153 12909 17187
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 13630 17144 13636 17196
rect 13688 17144 13694 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17153 15715 17187
rect 15856 17184 15884 17280
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15856 17156 15945 17184
rect 15657 17147 15715 17153
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 15672 17116 15700 17147
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 17589 17187 17647 17193
rect 17589 17184 17601 17187
rect 16632 17156 17601 17184
rect 16632 17144 16638 17156
rect 17589 17153 17601 17156
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 14056 17088 15976 17116
rect 14056 17076 14062 17088
rect 14936 17060 14964 17088
rect 5920 17020 6224 17048
rect 5813 17011 5871 17017
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 12621 17051 12679 17057
rect 12621 17048 12633 17051
rect 11112 17020 12633 17048
rect 11112 17008 11118 17020
rect 12621 17017 12633 17020
rect 12667 17017 12679 17051
rect 12621 17011 12679 17017
rect 14918 17008 14924 17060
rect 14976 17008 14982 17060
rect 15948 17048 15976 17088
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 16080 17088 18184 17116
rect 16080 17076 16086 17088
rect 16574 17048 16580 17060
rect 15212 17020 15884 17048
rect 15948 17020 16580 17048
rect 4948 16952 5028 16980
rect 4948 16940 4954 16952
rect 5074 16940 5080 16992
rect 5132 16940 5138 16992
rect 5902 16940 5908 16992
rect 5960 16980 5966 16992
rect 6914 16980 6920 16992
rect 5960 16952 6920 16980
rect 5960 16940 5966 16952
rect 6914 16940 6920 16952
rect 6972 16940 6978 16992
rect 8021 16983 8079 16989
rect 8021 16949 8033 16983
rect 8067 16980 8079 16983
rect 8110 16980 8116 16992
rect 8067 16952 8116 16980
rect 8067 16949 8079 16952
rect 8021 16943 8079 16949
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 15212 16980 15240 17020
rect 15856 16992 15884 17020
rect 16574 17008 16580 17020
rect 16632 17008 16638 17060
rect 18156 16992 18184 17088
rect 13596 16952 15240 16980
rect 13596 16940 13602 16952
rect 15378 16940 15384 16992
rect 15436 16940 15442 16992
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 17310 16980 17316 16992
rect 15896 16952 17316 16980
rect 15896 16940 15902 16952
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 18138 16940 18144 16992
rect 18196 16940 18202 16992
rect 1104 16890 19228 16912
rect 1104 16838 3215 16890
rect 3267 16838 3279 16890
rect 3331 16838 3343 16890
rect 3395 16838 3407 16890
rect 3459 16838 3471 16890
rect 3523 16838 7746 16890
rect 7798 16838 7810 16890
rect 7862 16838 7874 16890
rect 7926 16838 7938 16890
rect 7990 16838 8002 16890
rect 8054 16838 12277 16890
rect 12329 16838 12341 16890
rect 12393 16838 12405 16890
rect 12457 16838 12469 16890
rect 12521 16838 12533 16890
rect 12585 16838 16808 16890
rect 16860 16838 16872 16890
rect 16924 16838 16936 16890
rect 16988 16838 17000 16890
rect 17052 16838 17064 16890
rect 17116 16838 19228 16890
rect 1104 16816 19228 16838
rect 6454 16736 6460 16788
rect 6512 16776 6518 16788
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6512 16748 6561 16776
rect 6512 16736 6518 16748
rect 6549 16745 6561 16748
rect 6595 16745 6607 16779
rect 6549 16739 6607 16745
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8754 16776 8760 16788
rect 8536 16748 8760 16776
rect 8536 16736 8542 16748
rect 8754 16736 8760 16748
rect 8812 16776 8818 16788
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 8812 16748 8953 16776
rect 8812 16736 8818 16748
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10686 16776 10692 16788
rect 10192 16748 10692 16776
rect 10192 16736 10198 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 16758 16776 16764 16788
rect 15764 16748 16764 16776
rect 8110 16708 8116 16720
rect 7576 16680 8116 16708
rect 2866 16600 2872 16652
rect 2924 16600 2930 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4614 16640 4620 16652
rect 4111 16612 4620 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 7576 16649 7604 16680
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 8938 16640 8944 16652
rect 7699 16612 8944 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15764 16649 15792 16748
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 16022 16668 16028 16720
rect 16080 16668 16086 16720
rect 15749 16643 15807 16649
rect 15160 16612 15700 16640
rect 15160 16600 15166 16612
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3786 16572 3792 16584
rect 3191 16544 3792 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 2222 16464 2228 16516
rect 2280 16464 2286 16516
rect 3160 16504 3188 16535
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 5629 16575 5687 16581
rect 5629 16572 5641 16575
rect 5552 16544 5641 16572
rect 3068 16476 3188 16504
rect 3068 16448 3096 16476
rect 4522 16464 4528 16516
rect 4580 16464 4586 16516
rect 5552 16448 5580 16544
rect 5629 16541 5641 16544
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16541 6515 16575
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 6457 16535 6515 16541
rect 7668 16544 7757 16572
rect 6472 16448 6500 16535
rect 7668 16448 7696 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16572 7895 16575
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7883 16544 8125 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 8665 16575 8723 16581
rect 8665 16572 8677 16575
rect 8352 16544 8677 16572
rect 8352 16532 8358 16544
rect 8665 16541 8677 16544
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 15672 16572 15700 16612
rect 15749 16609 15761 16643
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 15838 16600 15844 16652
rect 15896 16600 15902 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16609 15991 16643
rect 15933 16603 15991 16609
rect 15948 16572 15976 16603
rect 16040 16581 16068 16668
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16640 16359 16643
rect 16666 16640 16672 16652
rect 16347 16612 16672 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16640 18107 16643
rect 18506 16640 18512 16652
rect 18095 16612 18512 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 18506 16600 18512 16612
rect 18564 16640 18570 16652
rect 18785 16643 18843 16649
rect 18785 16640 18797 16643
rect 18564 16612 18797 16640
rect 18564 16600 18570 16612
rect 18785 16609 18797 16612
rect 18831 16609 18843 16643
rect 18785 16603 18843 16609
rect 15672 16544 15976 16572
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 12158 16464 12164 16516
rect 12216 16464 12222 16516
rect 16577 16507 16635 16513
rect 16577 16473 16589 16507
rect 16623 16473 16635 16507
rect 16577 16467 16635 16473
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 2774 16436 2780 16448
rect 1443 16408 2780 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 2774 16396 2780 16408
rect 2832 16396 2838 16448
rect 3050 16396 3056 16448
rect 3108 16396 3114 16448
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 6270 16396 6276 16448
rect 6328 16396 6334 16448
rect 6454 16396 6460 16448
rect 6512 16396 6518 16448
rect 7374 16396 7380 16448
rect 7432 16396 7438 16448
rect 7650 16396 7656 16448
rect 7708 16396 7714 16448
rect 16209 16439 16267 16445
rect 16209 16405 16221 16439
rect 16255 16436 16267 16439
rect 16592 16436 16620 16467
rect 17310 16464 17316 16516
rect 17368 16464 17374 16516
rect 16255 16408 16620 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 18230 16396 18236 16448
rect 18288 16396 18294 16448
rect 1104 16346 19228 16368
rect 1104 16294 3875 16346
rect 3927 16294 3939 16346
rect 3991 16294 4003 16346
rect 4055 16294 4067 16346
rect 4119 16294 4131 16346
rect 4183 16294 8406 16346
rect 8458 16294 8470 16346
rect 8522 16294 8534 16346
rect 8586 16294 8598 16346
rect 8650 16294 8662 16346
rect 8714 16294 12937 16346
rect 12989 16294 13001 16346
rect 13053 16294 13065 16346
rect 13117 16294 13129 16346
rect 13181 16294 13193 16346
rect 13245 16294 17468 16346
rect 17520 16294 17532 16346
rect 17584 16294 17596 16346
rect 17648 16294 17660 16346
rect 17712 16294 17724 16346
rect 17776 16294 19228 16346
rect 1104 16272 19228 16294
rect 4522 16192 4528 16244
rect 4580 16192 4586 16244
rect 5534 16232 5540 16244
rect 5092 16204 5540 16232
rect 1578 16124 1584 16176
rect 1636 16164 1642 16176
rect 1857 16167 1915 16173
rect 1857 16164 1869 16167
rect 1636 16136 1869 16164
rect 1636 16124 1642 16136
rect 1857 16133 1869 16136
rect 1903 16133 1915 16167
rect 1857 16127 1915 16133
rect 5092 16105 5120 16204
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 6270 16192 6276 16244
rect 6328 16192 6334 16244
rect 8202 16192 8208 16244
rect 8260 16192 8266 16244
rect 8294 16192 8300 16244
rect 8352 16192 8358 16244
rect 8754 16192 8760 16244
rect 8812 16192 8818 16244
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9490 16232 9496 16244
rect 8987 16204 9496 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9732 16204 10456 16232
rect 9732 16192 9738 16204
rect 5258 16124 5264 16176
rect 5316 16164 5322 16176
rect 5353 16167 5411 16173
rect 5353 16164 5365 16167
rect 5316 16136 5365 16164
rect 5316 16124 5322 16136
rect 5353 16133 5365 16136
rect 5399 16133 5411 16167
rect 5353 16127 5411 16133
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 4632 15960 4660 16059
rect 5534 16056 5540 16108
rect 5592 16056 5598 16108
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16096 5779 16099
rect 6288 16096 6316 16192
rect 6822 16164 6828 16176
rect 6472 16136 6828 16164
rect 5767 16068 6316 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 6472 16105 6500 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 7466 16124 7472 16176
rect 7524 16124 7530 16176
rect 6457 16099 6515 16105
rect 6457 16096 6469 16099
rect 6420 16068 6469 16096
rect 6420 16056 6426 16068
rect 6457 16065 6469 16068
rect 6503 16065 6515 16099
rect 6457 16059 6515 16065
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5552 16028 5580 16056
rect 5215 16000 5580 16028
rect 6733 16031 6791 16037
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 6733 15997 6745 16031
rect 6779 16028 6791 16031
rect 7374 16028 7380 16040
rect 6779 16000 7380 16028
rect 6779 15997 6791 16000
rect 6733 15991 6791 15997
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8220 16028 8248 16192
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 8772 16096 8800 16192
rect 9858 16124 9864 16176
rect 9916 16124 9922 16176
rect 10428 16173 10456 16204
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 13265 16235 13323 16241
rect 13265 16232 13277 16235
rect 12860 16204 13277 16232
rect 12860 16192 12866 16204
rect 13265 16201 13277 16204
rect 13311 16201 13323 16235
rect 13265 16195 13323 16201
rect 16574 16192 16580 16244
rect 16632 16192 16638 16244
rect 16758 16192 16764 16244
rect 16816 16192 16822 16244
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 17368 16204 17417 16232
rect 17368 16192 17374 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 18230 16192 18236 16244
rect 18288 16192 18294 16244
rect 10413 16167 10471 16173
rect 10413 16133 10425 16167
rect 10459 16133 10471 16167
rect 10413 16127 10471 16133
rect 10704 16136 11560 16164
rect 10704 16108 10732 16136
rect 8527 16068 8800 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 10686 16056 10692 16108
rect 10744 16056 10750 16108
rect 11532 16105 11560 16136
rect 12066 16124 12072 16176
rect 12124 16164 12130 16176
rect 12124 16136 12282 16164
rect 12124 16124 12130 16136
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11517 16099 11575 16105
rect 11011 16068 11192 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 8220 16000 8677 16028
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 6454 15960 6460 15972
rect 4632 15932 6460 15960
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 11164 15904 11192 16068
rect 11517 16065 11529 16099
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11348 16000 11805 16028
rect 11348 15969 11376 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 13924 16028 13952 16059
rect 15654 16056 15660 16108
rect 15712 16056 15718 16108
rect 16592 16096 16620 16192
rect 16776 16164 16804 16192
rect 17681 16167 17739 16173
rect 17681 16164 17693 16167
rect 16776 16136 17693 16164
rect 17681 16133 17693 16136
rect 17727 16133 17739 16167
rect 17681 16127 17739 16133
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 16592 16068 17325 16096
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18248 16096 18276 16192
rect 18095 16068 18276 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 14918 16028 14924 16040
rect 13924 16000 14924 16028
rect 11793 15991 11851 15997
rect 14918 15988 14924 16000
rect 14976 15988 14982 16040
rect 17880 16028 17908 16059
rect 18506 16056 18512 16108
rect 18564 16056 18570 16108
rect 18601 16031 18659 16037
rect 18601 16028 18613 16031
rect 17880 16000 18613 16028
rect 18601 15997 18613 16000
rect 18647 16028 18659 16031
rect 18874 16028 18880 16040
rect 18647 16000 18880 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 18874 15988 18880 16000
rect 18932 15988 18938 16040
rect 11333 15963 11391 15969
rect 11333 15929 11345 15963
rect 11379 15929 11391 15963
rect 11333 15923 11391 15929
rect 18138 15920 18144 15972
rect 18196 15920 18202 15972
rect 2133 15895 2191 15901
rect 2133 15861 2145 15895
rect 2179 15892 2191 15895
rect 4246 15892 4252 15904
rect 2179 15864 4252 15892
rect 2179 15861 2191 15864
rect 2133 15855 2191 15861
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 5074 15892 5080 15904
rect 4755 15864 5080 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 11146 15852 11152 15904
rect 11204 15852 11210 15904
rect 13814 15852 13820 15904
rect 13872 15852 13878 15904
rect 15565 15895 15623 15901
rect 15565 15861 15577 15895
rect 15611 15892 15623 15895
rect 16114 15892 16120 15904
rect 15611 15864 16120 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 1104 15802 19228 15824
rect 1104 15750 3215 15802
rect 3267 15750 3279 15802
rect 3331 15750 3343 15802
rect 3395 15750 3407 15802
rect 3459 15750 3471 15802
rect 3523 15750 7746 15802
rect 7798 15750 7810 15802
rect 7862 15750 7874 15802
rect 7926 15750 7938 15802
rect 7990 15750 8002 15802
rect 8054 15750 12277 15802
rect 12329 15750 12341 15802
rect 12393 15750 12405 15802
rect 12457 15750 12469 15802
rect 12521 15750 12533 15802
rect 12585 15750 16808 15802
rect 16860 15750 16872 15802
rect 16924 15750 16936 15802
rect 16988 15750 17000 15802
rect 17052 15750 17064 15802
rect 17116 15750 19228 15802
rect 1104 15728 19228 15750
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7466 15688 7472 15700
rect 7423 15660 7472 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 9858 15648 9864 15700
rect 9916 15648 9922 15700
rect 11146 15648 11152 15700
rect 11204 15648 11210 15700
rect 11977 15691 12035 15697
rect 11977 15657 11989 15691
rect 12023 15688 12035 15691
rect 12066 15688 12072 15700
rect 12023 15660 12072 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 13814 15648 13820 15700
rect 13872 15648 13878 15700
rect 8110 15620 8116 15632
rect 8036 15592 8116 15620
rect 2222 15512 2228 15564
rect 2280 15512 2286 15564
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15552 2743 15555
rect 2774 15552 2780 15564
rect 2731 15524 2780 15552
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 2774 15512 2780 15524
rect 2832 15552 2838 15564
rect 3418 15552 3424 15564
rect 2832 15524 3424 15552
rect 2832 15512 2838 15524
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 8036 15561 8064 15592
rect 8110 15580 8116 15592
rect 8168 15580 8174 15632
rect 8481 15623 8539 15629
rect 8481 15589 8493 15623
rect 8527 15620 8539 15623
rect 8754 15620 8760 15632
rect 8527 15592 8760 15620
rect 8527 15589 8539 15592
rect 8481 15583 8539 15589
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10962 15620 10968 15632
rect 10008 15592 10968 15620
rect 10008 15580 10014 15592
rect 10962 15580 10968 15592
rect 11020 15620 11026 15632
rect 11020 15592 11928 15620
rect 11020 15580 11026 15592
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15521 8079 15555
rect 8665 15555 8723 15561
rect 8665 15552 8677 15555
rect 8021 15515 8079 15521
rect 8128 15524 8677 15552
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 3142 15484 3148 15496
rect 2639 15456 3148 15484
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 3142 15444 3148 15456
rect 3200 15484 3206 15496
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 3200 15456 4353 15484
rect 3200 15444 3206 15456
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 6454 15484 6460 15496
rect 4341 15447 4399 15453
rect 6288 15456 6460 15484
rect 6288 15360 6316 15456
rect 6454 15444 6460 15456
rect 6512 15484 6518 15496
rect 8128 15493 8156 15524
rect 8665 15521 8677 15524
rect 8711 15521 8723 15555
rect 8665 15515 8723 15521
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 6512 15456 7297 15484
rect 6512 15444 6518 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7285 15447 7343 15453
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 8938 15484 8944 15496
rect 8803 15456 8944 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 8588 15416 8616 15447
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9968 15493 9996 15580
rect 10778 15512 10784 15564
rect 10836 15512 10842 15564
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 10796 15484 10824 15512
rect 11900 15493 11928 15592
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15552 12219 15555
rect 13630 15552 13636 15564
rect 12207 15524 13636 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10796 15456 11069 15484
rect 9953 15447 10011 15453
rect 11057 15453 11069 15456
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11885 15487 11943 15493
rect 11287 15456 11560 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 6972 15388 8616 15416
rect 6972 15376 6978 15388
rect 11532 15360 11560 15456
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 13832 15484 13860 15648
rect 13909 15555 13967 15561
rect 13909 15521 13921 15555
rect 13955 15552 13967 15555
rect 14458 15552 14464 15564
rect 13955 15524 14464 15552
rect 13955 15521 13967 15524
rect 13909 15515 13967 15521
rect 14458 15512 14464 15524
rect 14516 15552 14522 15564
rect 14553 15555 14611 15561
rect 14553 15552 14565 15555
rect 14516 15524 14565 15552
rect 14516 15512 14522 15524
rect 14553 15521 14565 15524
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15552 15255 15555
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15243 15524 15669 15552
rect 15243 15521 15255 15524
rect 15197 15515 15255 15521
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 13570 15456 13860 15484
rect 11885 15447 11943 15453
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15436 15456 15485 15484
rect 15436 15444 15442 15456
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 12434 15376 12440 15428
rect 12492 15376 12498 15428
rect 3786 15308 3792 15360
rect 3844 15308 3850 15360
rect 6270 15308 6276 15360
rect 6328 15308 6334 15360
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 13906 15348 13912 15360
rect 11572 15320 13912 15348
rect 11572 15308 11578 15320
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 14274 15308 14280 15360
rect 14332 15348 14338 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 14332 15320 15301 15348
rect 14332 15308 14338 15320
rect 15289 15317 15301 15320
rect 15335 15317 15347 15351
rect 15289 15311 15347 15317
rect 1104 15258 19228 15280
rect 1104 15206 3875 15258
rect 3927 15206 3939 15258
rect 3991 15206 4003 15258
rect 4055 15206 4067 15258
rect 4119 15206 4131 15258
rect 4183 15206 8406 15258
rect 8458 15206 8470 15258
rect 8522 15206 8534 15258
rect 8586 15206 8598 15258
rect 8650 15206 8662 15258
rect 8714 15206 12937 15258
rect 12989 15206 13001 15258
rect 13053 15206 13065 15258
rect 13117 15206 13129 15258
rect 13181 15206 13193 15258
rect 13245 15206 17468 15258
rect 17520 15206 17532 15258
rect 17584 15206 17596 15258
rect 17648 15206 17660 15258
rect 17712 15206 17724 15258
rect 17776 15206 19228 15258
rect 1104 15184 19228 15206
rect 3142 15104 3148 15156
rect 3200 15104 3206 15156
rect 7190 15104 7196 15156
rect 7248 15104 7254 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12492 15116 13093 15144
rect 12492 15104 12498 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 13446 15104 13452 15156
rect 13504 15104 13510 15156
rect 15746 15104 15752 15156
rect 15804 15104 15810 15156
rect 2130 15036 2136 15088
rect 2188 15036 2194 15088
rect 7101 15079 7159 15085
rect 7101 15076 7113 15079
rect 6748 15048 7113 15076
rect 3418 14968 3424 15020
rect 3476 14968 3482 15020
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3786 15008 3792 15020
rect 3651 14980 3792 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 6748 15017 6776 15048
rect 7101 15045 7113 15048
rect 7147 15045 7159 15079
rect 7101 15039 7159 15045
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7208 15017 7236 15104
rect 10410 15076 10416 15088
rect 9876 15048 10416 15076
rect 7009 15011 7067 15017
rect 7009 15008 7021 15011
rect 6972 14980 7021 15008
rect 6972 14968 6978 14980
rect 7009 14977 7021 14980
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 9876 14952 9904 15048
rect 10410 15036 10416 15048
rect 10468 15076 10474 15088
rect 10468 15048 10916 15076
rect 10468 15036 10474 15048
rect 10778 14968 10784 15020
rect 10836 14968 10842 15020
rect 10888 15017 10916 15048
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 13464 15008 13492 15104
rect 15764 15076 15792 15104
rect 14200 15048 15516 15076
rect 15764 15048 16160 15076
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 13403 14980 13737 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 13725 14977 13737 14980
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 14200 15008 14228 15048
rect 13964 14980 14228 15008
rect 13964 14968 13970 14980
rect 14274 14968 14280 15020
rect 14332 14968 14338 15020
rect 14458 14968 14464 15020
rect 14516 14968 14522 15020
rect 1394 14900 1400 14952
rect 1452 14900 1458 14952
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 6871 14912 7052 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 2832 14844 3249 14872
rect 2832 14832 2838 14844
rect 3237 14841 3249 14844
rect 3283 14841 3295 14875
rect 3237 14835 3295 14841
rect 7024 14816 7052 14912
rect 9858 14900 9864 14952
rect 9916 14900 9922 14952
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11011 14912 11529 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 10704 14872 10732 14903
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 11756 14912 12081 14940
rect 11756 14900 11762 14912
rect 12069 14909 12081 14912
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 13265 14943 13323 14949
rect 13265 14909 13277 14943
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13280 14872 13308 14903
rect 13446 14900 13452 14952
rect 13504 14900 13510 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 14292 14940 14320 14968
rect 13587 14912 14320 14940
rect 14553 14943 14611 14949
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 15378 14940 15384 14952
rect 14599 14912 15384 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15488 14940 15516 15048
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 15008 15899 15011
rect 16022 15008 16028 15020
rect 15887 14980 16028 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16132 15017 16160 15048
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16316 14940 16344 14971
rect 17494 14968 17500 15020
rect 17552 14968 17558 15020
rect 15488 14912 16344 14940
rect 17589 14943 17647 14949
rect 16132 14884 16160 14912
rect 17589 14909 17601 14943
rect 17635 14940 17647 14943
rect 18230 14940 18236 14952
rect 17635 14912 18236 14940
rect 17635 14909 17647 14912
rect 17589 14903 17647 14909
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 14093 14875 14151 14881
rect 14093 14872 14105 14875
rect 10704 14844 10916 14872
rect 13280 14844 14105 14872
rect 10888 14816 10916 14844
rect 13556 14816 13584 14844
rect 14093 14841 14105 14844
rect 14139 14841 14151 14875
rect 14093 14835 14151 14841
rect 16114 14832 16120 14884
rect 16172 14832 16178 14884
rect 6454 14764 6460 14816
rect 6512 14764 6518 14816
rect 7006 14764 7012 14816
rect 7064 14764 7070 14816
rect 10502 14764 10508 14816
rect 10560 14764 10566 14816
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 13538 14764 13544 14816
rect 13596 14764 13602 14816
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 15930 14764 15936 14816
rect 15988 14764 15994 14816
rect 16209 14807 16267 14813
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 16574 14804 16580 14816
rect 16255 14776 16580 14804
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 17862 14804 17868 14816
rect 17175 14776 17868 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 1104 14714 19228 14736
rect 1104 14662 3215 14714
rect 3267 14662 3279 14714
rect 3331 14662 3343 14714
rect 3395 14662 3407 14714
rect 3459 14662 3471 14714
rect 3523 14662 7746 14714
rect 7798 14662 7810 14714
rect 7862 14662 7874 14714
rect 7926 14662 7938 14714
rect 7990 14662 8002 14714
rect 8054 14662 12277 14714
rect 12329 14662 12341 14714
rect 12393 14662 12405 14714
rect 12457 14662 12469 14714
rect 12521 14662 12533 14714
rect 12585 14662 16808 14714
rect 16860 14662 16872 14714
rect 16924 14662 16936 14714
rect 16988 14662 17000 14714
rect 17052 14662 17064 14714
rect 17116 14662 19228 14714
rect 1104 14640 19228 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2317 14603 2375 14609
rect 2317 14600 2329 14603
rect 1728 14572 2329 14600
rect 1728 14560 1734 14572
rect 2317 14569 2329 14572
rect 2363 14569 2375 14603
rect 2317 14563 2375 14569
rect 5534 14560 5540 14612
rect 5592 14560 5598 14612
rect 6454 14560 6460 14612
rect 6512 14560 6518 14612
rect 7006 14560 7012 14612
rect 7064 14560 7070 14612
rect 9858 14560 9864 14612
rect 9916 14560 9922 14612
rect 10124 14603 10182 14609
rect 10124 14569 10136 14603
rect 10170 14600 10182 14603
rect 10502 14600 10508 14612
rect 10170 14572 10508 14600
rect 10170 14569 10182 14572
rect 10124 14563 10182 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 12529 14603 12587 14609
rect 12529 14600 12541 14603
rect 10928 14572 12541 14600
rect 10928 14560 10934 14572
rect 12529 14569 12541 14572
rect 12575 14569 12587 14603
rect 13538 14600 13544 14612
rect 12529 14563 12587 14569
rect 13464 14572 13544 14600
rect 2130 14492 2136 14544
rect 2188 14492 2194 14544
rect 2222 14424 2228 14476
rect 2280 14464 2286 14476
rect 2501 14467 2559 14473
rect 2501 14464 2513 14467
rect 2280 14436 2513 14464
rect 2280 14424 2286 14436
rect 2501 14433 2513 14436
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 2774 14424 2780 14476
rect 2832 14424 2838 14476
rect 3050 14424 3056 14476
rect 3108 14464 3114 14476
rect 4065 14467 4123 14473
rect 3108 14436 3832 14464
rect 3108 14424 3114 14436
rect 3804 14408 3832 14436
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 6472 14464 6500 14560
rect 6730 14492 6736 14544
rect 6788 14532 6794 14544
rect 7650 14532 7656 14544
rect 6788 14504 7656 14532
rect 6788 14492 6794 14504
rect 7650 14492 7656 14504
rect 7708 14532 7714 14544
rect 9876 14532 9904 14560
rect 7708 14504 9904 14532
rect 7708 14492 7714 14504
rect 4111 14436 6500 14464
rect 6549 14467 6607 14473
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 7098 14464 7104 14476
rect 6595 14436 7104 14464
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 7098 14424 7104 14436
rect 7156 14464 7162 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7156 14436 7573 14464
rect 7156 14424 7162 14436
rect 7561 14433 7573 14436
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14464 9919 14467
rect 10686 14464 10692 14476
rect 9907 14436 10692 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 11655 14436 12357 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 12345 14433 12357 14436
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 2038 14356 2044 14408
rect 2096 14356 2102 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 2608 14328 2636 14359
rect 2682 14356 2688 14408
rect 2740 14356 2746 14408
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14396 3203 14399
rect 3191 14368 3740 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 2976 14328 3004 14359
rect 3712 14340 3740 14368
rect 3786 14356 3792 14408
rect 3844 14356 3850 14408
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 2608 14300 3188 14328
rect 3050 14220 3056 14272
rect 3108 14220 3114 14272
rect 3160 14260 3188 14300
rect 3694 14288 3700 14340
rect 3752 14288 3758 14340
rect 5721 14331 5779 14337
rect 5721 14328 5733 14331
rect 5290 14300 5733 14328
rect 5721 14297 5733 14300
rect 5767 14297 5779 14331
rect 5828 14328 5856 14359
rect 6270 14328 6276 14340
rect 5828 14300 6276 14328
rect 5721 14291 5779 14297
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 6656 14328 6684 14359
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7466 14396 7472 14408
rect 6871 14368 7472 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14365 9091 14399
rect 12360 14396 12388 14427
rect 12802 14424 12808 14476
rect 12860 14424 12866 14476
rect 13464 14473 13492 14572
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13814 14560 13820 14612
rect 13872 14560 13878 14612
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 16942 14600 16948 14612
rect 16807 14572 16948 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 16942 14560 16948 14572
rect 17000 14600 17006 14612
rect 17494 14600 17500 14612
rect 17000 14572 17500 14600
rect 17000 14560 17006 14572
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 18874 14560 18880 14612
rect 18932 14560 18938 14612
rect 13832 14532 13860 14560
rect 13556 14504 13860 14532
rect 13449 14467 13507 14473
rect 13449 14433 13461 14467
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 13556 14405 13584 14504
rect 13630 14424 13636 14476
rect 13688 14464 13694 14476
rect 14366 14464 14372 14476
rect 13688 14436 14372 14464
rect 13688 14424 13694 14436
rect 14366 14424 14372 14436
rect 14424 14464 14430 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14424 14436 15025 14464
rect 14424 14424 14430 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 16724 14436 17141 14464
rect 16724 14424 16730 14436
rect 17129 14433 17141 14436
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 12897 14399 12955 14405
rect 12897 14396 12909 14399
rect 12360 14368 12909 14396
rect 9033 14359 9091 14365
rect 12897 14365 12909 14368
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 7190 14328 7196 14340
rect 6656 14300 7196 14328
rect 7190 14288 7196 14300
rect 7248 14288 7254 14340
rect 9048 14272 9076 14359
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 10870 14288 10876 14340
rect 10928 14288 10934 14340
rect 15286 14288 15292 14340
rect 15344 14288 15350 14340
rect 15930 14288 15936 14340
rect 15988 14288 15994 14340
rect 17310 14288 17316 14340
rect 17368 14328 17374 14340
rect 17405 14331 17463 14337
rect 17405 14328 17417 14331
rect 17368 14300 17417 14328
rect 17368 14288 17374 14300
rect 17405 14297 17417 14300
rect 17451 14297 17463 14331
rect 17405 14291 17463 14297
rect 4982 14260 4988 14272
rect 3160 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 6365 14263 6423 14269
rect 6365 14229 6377 14263
rect 6411 14260 6423 14263
rect 6546 14260 6552 14272
rect 6411 14232 6552 14260
rect 6411 14229 6423 14232
rect 6365 14223 6423 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 9030 14220 9036 14272
rect 9088 14220 9094 14272
rect 9122 14220 9128 14272
rect 9180 14220 9186 14272
rect 11790 14220 11796 14272
rect 11848 14220 11854 14272
rect 13173 14263 13231 14269
rect 13173 14229 13185 14263
rect 13219 14260 13231 14263
rect 13262 14260 13268 14272
rect 13219 14232 13268 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 16022 14220 16028 14272
rect 16080 14260 16086 14272
rect 16298 14260 16304 14272
rect 16080 14232 16304 14260
rect 16080 14220 16086 14232
rect 16298 14220 16304 14232
rect 16356 14260 16362 14272
rect 18046 14260 18052 14272
rect 16356 14232 18052 14260
rect 16356 14220 16362 14232
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 1104 14170 19228 14192
rect 1104 14118 3875 14170
rect 3927 14118 3939 14170
rect 3991 14118 4003 14170
rect 4055 14118 4067 14170
rect 4119 14118 4131 14170
rect 4183 14118 8406 14170
rect 8458 14118 8470 14170
rect 8522 14118 8534 14170
rect 8586 14118 8598 14170
rect 8650 14118 8662 14170
rect 8714 14118 12937 14170
rect 12989 14118 13001 14170
rect 13053 14118 13065 14170
rect 13117 14118 13129 14170
rect 13181 14118 13193 14170
rect 13245 14118 17468 14170
rect 17520 14118 17532 14170
rect 17584 14118 17596 14170
rect 17648 14118 17660 14170
rect 17712 14118 17724 14170
rect 17776 14118 19228 14170
rect 1104 14096 19228 14118
rect 3050 14056 3056 14068
rect 2746 14028 3056 14056
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 2746 13920 2774 14028
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 6089 14059 6147 14065
rect 6089 14025 6101 14059
rect 6135 14056 6147 14059
rect 6135 14028 6960 14056
rect 6135 14025 6147 14028
rect 6089 14019 6147 14025
rect 4246 13948 4252 14000
rect 4304 13988 4310 14000
rect 4617 13991 4675 13997
rect 4617 13988 4629 13991
rect 4304 13960 4629 13988
rect 4304 13948 4310 13960
rect 4617 13957 4629 13960
rect 4663 13988 4675 13991
rect 4890 13988 4896 14000
rect 4663 13960 4896 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 6546 13948 6552 14000
rect 6604 13988 6610 14000
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 6604 13960 6653 13988
rect 6604 13948 6610 13960
rect 6641 13957 6653 13960
rect 6687 13957 6699 13991
rect 6932 13988 6960 14028
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 10965 14059 11023 14065
rect 10965 14056 10977 14059
rect 10928 14028 10977 14056
rect 10928 14016 10934 14028
rect 10965 14025 10977 14028
rect 11011 14025 11023 14059
rect 10965 14019 11023 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11698 14056 11704 14068
rect 11563 14028 11704 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11790 14016 11796 14068
rect 11848 14016 11854 14068
rect 13538 14016 13544 14068
rect 13596 14016 13602 14068
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 15344 14028 15669 14056
rect 15344 14016 15350 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 18506 14016 18512 14068
rect 18564 14016 18570 14068
rect 6932 13960 7130 13988
rect 6641 13951 6699 13957
rect 9122 13948 9128 14000
rect 9180 13948 9186 14000
rect 2455 13892 2774 13920
rect 5997 13923 6055 13929
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 5997 13889 6009 13923
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 2280 13824 2329 13852
rect 2280 13812 2286 13824
rect 2317 13821 2329 13824
rect 2363 13821 2375 13855
rect 6012 13852 6040 13883
rect 8294 13880 8300 13932
rect 8352 13880 8358 13932
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 10962 13920 10968 13932
rect 10919 13892 10968 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11808 13929 11836 14016
rect 13556 13988 13584 14016
rect 14829 13991 14887 13997
rect 14829 13988 14841 13991
rect 12912 13960 13584 13988
rect 14398 13960 14841 13988
rect 12912 13929 12940 13960
rect 14829 13957 14841 13960
rect 14875 13957 14887 13991
rect 17862 13988 17868 14000
rect 14829 13951 14887 13957
rect 15856 13960 17868 13988
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 6270 13852 6276 13864
rect 6012 13824 6276 13852
rect 2317 13815 2375 13821
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 6362 13812 6368 13864
rect 6420 13812 6426 13864
rect 11716 13852 11744 13883
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 15746 13880 15752 13932
rect 15804 13880 15810 13932
rect 15856 13929 15884 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 18064 13988 18092 14016
rect 18064 13960 18460 13988
rect 15841 13923 15899 13929
rect 15841 13889 15853 13923
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 16163 13892 17969 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13920 18199 13923
rect 18230 13920 18236 13932
rect 18187 13892 18236 13920
rect 18187 13889 18199 13892
rect 18141 13883 18199 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18432 13929 18460 13960
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 12802 13852 12808 13864
rect 11716 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13262 13852 13268 13864
rect 13219 13824 13268 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 14642 13812 14648 13864
rect 14700 13812 14706 13864
rect 15764 13852 15792 13880
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15764 13824 15945 13852
rect 15933 13821 15945 13824
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13821 16083 13855
rect 16025 13815 16083 13821
rect 3694 13744 3700 13796
rect 3752 13784 3758 13796
rect 3752 13756 4936 13784
rect 3752 13744 3758 13756
rect 2685 13719 2743 13725
rect 2685 13685 2697 13719
rect 2731 13716 2743 13719
rect 4246 13716 4252 13728
rect 2731 13688 4252 13716
rect 2731 13685 2743 13688
rect 2685 13679 2743 13685
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 4908 13725 4936 13756
rect 15654 13744 15660 13796
rect 15712 13784 15718 13796
rect 15838 13784 15844 13796
rect 15712 13756 15844 13784
rect 15712 13744 15718 13756
rect 15838 13744 15844 13756
rect 15896 13784 15902 13796
rect 16040 13784 16068 13815
rect 16942 13812 16948 13864
rect 17000 13852 17006 13864
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 17000 13824 17233 13852
rect 17000 13812 17006 13824
rect 17221 13821 17233 13824
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 17865 13855 17923 13861
rect 17865 13821 17877 13855
rect 17911 13852 17923 13855
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 17911 13824 18337 13852
rect 17911 13821 17923 13824
rect 17865 13815 17923 13821
rect 18325 13821 18337 13824
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 15896 13756 16068 13784
rect 15896 13744 15902 13756
rect 4893 13719 4951 13725
rect 4893 13685 4905 13719
rect 4939 13716 4951 13719
rect 7006 13716 7012 13728
rect 4939 13688 7012 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 8110 13676 8116 13728
rect 8168 13676 8174 13728
rect 8560 13719 8618 13725
rect 8560 13685 8572 13719
rect 8606 13716 8618 13719
rect 8754 13716 8760 13728
rect 8606 13688 8760 13716
rect 8606 13685 8618 13688
rect 8560 13679 8618 13685
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 10042 13676 10048 13728
rect 10100 13676 10106 13728
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 17218 13716 17224 13728
rect 17092 13688 17224 13716
rect 17092 13676 17098 13688
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 1104 13626 19228 13648
rect 1104 13574 3215 13626
rect 3267 13574 3279 13626
rect 3331 13574 3343 13626
rect 3395 13574 3407 13626
rect 3459 13574 3471 13626
rect 3523 13574 7746 13626
rect 7798 13574 7810 13626
rect 7862 13574 7874 13626
rect 7926 13574 7938 13626
rect 7990 13574 8002 13626
rect 8054 13574 12277 13626
rect 12329 13574 12341 13626
rect 12393 13574 12405 13626
rect 12457 13574 12469 13626
rect 12521 13574 12533 13626
rect 12585 13574 16808 13626
rect 16860 13574 16872 13626
rect 16924 13574 16936 13626
rect 16988 13574 17000 13626
rect 17052 13574 17064 13626
rect 17116 13574 19228 13626
rect 1104 13552 19228 13574
rect 6362 13472 6368 13524
rect 6420 13512 6426 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 6420 13484 6561 13512
rect 6420 13472 6426 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 6549 13475 6607 13481
rect 7098 13472 7104 13524
rect 7156 13472 7162 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 12802 13512 12808 13524
rect 12575 13484 12808 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 17129 13515 17187 13521
rect 17129 13481 17141 13515
rect 17175 13512 17187 13515
rect 17310 13512 17316 13524
rect 17175 13484 17316 13512
rect 17175 13481 17187 13484
rect 17129 13475 17187 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 7650 13444 7656 13456
rect 7392 13416 7656 13444
rect 4614 13336 4620 13388
rect 4672 13336 4678 13388
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 6178 13376 6184 13388
rect 5123 13348 6184 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 7392 13385 7420 13416
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13345 7435 13379
rect 8110 13376 8116 13388
rect 7377 13339 7435 13345
rect 7484 13348 8116 13376
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 2096 13280 3801 13308
rect 2096 13268 2102 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5626 13308 5632 13320
rect 5031 13280 5632 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 7484 13317 7512 13348
rect 8110 13336 8116 13348
rect 8168 13376 8174 13388
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 8168 13348 8677 13376
rect 8168 13336 8174 13348
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 10686 13336 10692 13388
rect 10744 13376 10750 13388
rect 10781 13379 10839 13385
rect 10781 13376 10793 13379
rect 10744 13348 10793 13376
rect 10744 13336 10750 13348
rect 10781 13345 10793 13348
rect 10827 13345 10839 13379
rect 10781 13339 10839 13345
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13376 17003 13379
rect 17862 13376 17868 13388
rect 16991 13348 17868 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13308 8999 13311
rect 9030 13308 9036 13320
rect 8987 13280 9036 13308
rect 8987 13277 8999 13280
rect 8941 13271 8999 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13308 9643 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9631 13280 9689 13308
rect 9631 13277 9643 13280
rect 9585 13271 9643 13277
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 5258 13200 5264 13252
rect 5316 13200 5322 13252
rect 9416 13240 9444 13271
rect 10042 13268 10048 13320
rect 10100 13268 10106 13320
rect 10226 13268 10232 13320
rect 10284 13268 10290 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 16632 13280 16865 13308
rect 16632 13268 16638 13280
rect 16853 13277 16865 13280
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 10060 13240 10088 13268
rect 9416 13212 10088 13240
rect 11054 13200 11060 13252
rect 11112 13200 11118 13252
rect 11790 13200 11796 13252
rect 11848 13200 11854 13252
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4890 13172 4896 13184
rect 3927 13144 4896 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 8110 13132 8116 13184
rect 8168 13132 8174 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8996 13144 9045 13172
rect 8996 13132 9002 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 9214 13132 9220 13184
rect 9272 13132 9278 13184
rect 1104 13082 19228 13104
rect 1104 13030 3875 13082
rect 3927 13030 3939 13082
rect 3991 13030 4003 13082
rect 4055 13030 4067 13082
rect 4119 13030 4131 13082
rect 4183 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 8534 13082
rect 8586 13030 8598 13082
rect 8650 13030 8662 13082
rect 8714 13030 12937 13082
rect 12989 13030 13001 13082
rect 13053 13030 13065 13082
rect 13117 13030 13129 13082
rect 13181 13030 13193 13082
rect 13245 13030 17468 13082
rect 17520 13030 17532 13082
rect 17584 13030 17596 13082
rect 17648 13030 17660 13082
rect 17712 13030 17724 13082
rect 17776 13030 19228 13082
rect 1104 13008 19228 13030
rect 4890 12928 4896 12980
rect 4948 12928 4954 12980
rect 6178 12928 6184 12980
rect 6236 12928 6242 12980
rect 7466 12928 7472 12980
rect 7524 12928 7530 12980
rect 8110 12968 8116 12980
rect 7852 12940 8116 12968
rect 4246 12860 4252 12912
rect 4304 12900 4310 12912
rect 4709 12903 4767 12909
rect 4709 12900 4721 12903
rect 4304 12872 4721 12900
rect 4304 12860 4310 12872
rect 4709 12869 4721 12872
rect 4755 12869 4767 12903
rect 4908 12900 4936 12928
rect 4908 12872 5198 12900
rect 4709 12863 4767 12869
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2682 12832 2688 12844
rect 2639 12804 2688 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 7650 12792 7656 12844
rect 7708 12792 7714 12844
rect 7852 12841 7880 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 9677 12971 9735 12977
rect 9677 12937 9689 12971
rect 9723 12968 9735 12971
rect 10226 12968 10232 12980
rect 9723 12940 10232 12968
rect 9723 12937 9735 12940
rect 9677 12931 9735 12937
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 11054 12928 11060 12980
rect 11112 12928 11118 12980
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 11790 12928 11796 12980
rect 11848 12928 11854 12980
rect 14277 12971 14335 12977
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 14366 12968 14372 12980
rect 14323 12940 14372 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 18230 12928 18236 12980
rect 18288 12968 18294 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 18288 12940 18889 12968
rect 18288 12928 18294 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 8294 12900 8300 12912
rect 7944 12872 8300 12900
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 7944 12773 7972 12872
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 8938 12860 8944 12912
rect 8996 12860 9002 12912
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10244 12832 10272 12928
rect 11164 12900 11192 12928
rect 11164 12872 11744 12900
rect 10183 12804 10272 12832
rect 10689 12835 10747 12841
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 11238 12832 11244 12844
rect 10735 12804 11244 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11716 12841 11744 12872
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 12676 12872 13001 12900
rect 12676 12860 12682 12872
rect 12989 12869 13001 12872
rect 13035 12869 13047 12903
rect 12989 12863 13047 12869
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 15488 12832 15516 12928
rect 18414 12860 18420 12912
rect 18472 12860 18478 12912
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 15488 12804 15577 12832
rect 11701 12795 11759 12801
rect 15565 12801 15577 12804
rect 15611 12832 15623 12835
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15611 12804 15945 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 15933 12801 15945 12804
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 16724 12804 17141 12832
rect 16724 12792 16730 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 3896 12736 4445 12764
rect 3896 12640 3924 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12764 8263 12767
rect 8938 12764 8944 12776
rect 8251 12736 8944 12764
rect 8251 12733 8263 12736
rect 8205 12727 8263 12733
rect 6362 12656 6368 12708
rect 6420 12696 6426 12708
rect 7944 12696 7972 12727
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 10042 12724 10048 12776
rect 10100 12724 10106 12776
rect 10594 12724 10600 12776
rect 10652 12724 10658 12776
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 6420 12668 7972 12696
rect 15488 12696 15516 12727
rect 15654 12724 15660 12776
rect 15712 12724 15718 12776
rect 15746 12724 15752 12776
rect 15804 12724 15810 12776
rect 17402 12724 17408 12776
rect 17460 12724 17466 12776
rect 16666 12696 16672 12708
rect 15488 12668 16672 12696
rect 6420 12656 6426 12668
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 3878 12588 3884 12640
rect 3936 12588 3942 12640
rect 9766 12588 9772 12640
rect 9824 12588 9830 12640
rect 15286 12588 15292 12640
rect 15344 12588 15350 12640
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 18046 12628 18052 12640
rect 16071 12600 18052 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 1104 12538 19228 12560
rect 1104 12486 3215 12538
rect 3267 12486 3279 12538
rect 3331 12486 3343 12538
rect 3395 12486 3407 12538
rect 3459 12486 3471 12538
rect 3523 12486 7746 12538
rect 7798 12486 7810 12538
rect 7862 12486 7874 12538
rect 7926 12486 7938 12538
rect 7990 12486 8002 12538
rect 8054 12486 12277 12538
rect 12329 12486 12341 12538
rect 12393 12486 12405 12538
rect 12457 12486 12469 12538
rect 12521 12486 12533 12538
rect 12585 12486 16808 12538
rect 16860 12486 16872 12538
rect 16924 12486 16936 12538
rect 16988 12486 17000 12538
rect 17052 12486 17064 12538
rect 17116 12486 19228 12538
rect 1104 12464 19228 12486
rect 5626 12384 5632 12436
rect 5684 12384 5690 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7708 12396 7849 12424
rect 7708 12384 7714 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12393 9827 12427
rect 9769 12387 9827 12393
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 3878 12288 3884 12300
rect 1452 12260 3884 12288
rect 1452 12248 1458 12260
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 5644 12288 5672 12384
rect 5994 12316 6000 12368
rect 6052 12356 6058 12368
rect 6270 12356 6276 12368
rect 6052 12328 6276 12356
rect 6052 12316 6058 12328
rect 6270 12316 6276 12328
rect 6328 12356 6334 12368
rect 9030 12356 9036 12368
rect 6328 12328 9036 12356
rect 6328 12316 6334 12328
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5644 12260 5733 12288
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 6454 12180 6460 12232
rect 6512 12180 6518 12232
rect 6840 12229 6868 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 9784 12300 9812 12387
rect 11238 12384 11244 12436
rect 11296 12384 11302 12436
rect 18414 12384 18420 12436
rect 18472 12384 18478 12436
rect 17402 12316 17408 12368
rect 17460 12356 17466 12368
rect 17681 12359 17739 12365
rect 17681 12356 17693 12359
rect 17460 12328 17693 12356
rect 17460 12316 17466 12328
rect 17681 12325 17693 12328
rect 17727 12325 17739 12359
rect 17681 12319 17739 12325
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 14553 12291 14611 12297
rect 13004 12260 13768 12288
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8168 12192 8401 12220
rect 8168 12180 8174 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11514 12220 11520 12232
rect 11379 12192 11520 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 1670 12112 1676 12164
rect 1728 12112 1734 12164
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 4157 12155 4215 12161
rect 2004 12124 2162 12152
rect 2004 12112 2010 12124
rect 4157 12121 4169 12155
rect 4203 12152 4215 12155
rect 4246 12152 4252 12164
rect 4203 12124 4252 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 6549 12155 6607 12161
rect 6549 12152 6561 12155
rect 5382 12124 6561 12152
rect 6549 12121 6561 12124
rect 6595 12121 6607 12155
rect 6549 12115 6607 12121
rect 11054 12112 11060 12164
rect 11112 12112 11118 12164
rect 11164 12152 11192 12183
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 13004 12229 13032 12260
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 13219 12192 13308 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 11422 12152 11428 12164
rect 11164 12124 11428 12152
rect 11164 12096 11192 12124
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 3016 12056 3157 12084
rect 3016 12044 3022 12056
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3145 12047 3203 12053
rect 6270 12044 6276 12096
rect 6328 12084 6334 12096
rect 6365 12087 6423 12093
rect 6365 12084 6377 12087
rect 6328 12056 6377 12084
rect 6328 12044 6334 12056
rect 6365 12053 6377 12056
rect 6411 12053 6423 12087
rect 6365 12047 6423 12053
rect 6914 12044 6920 12096
rect 6972 12044 6978 12096
rect 11146 12044 11152 12096
rect 11204 12044 11210 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 13280 12093 13308 12192
rect 13740 12152 13768 12260
rect 14553 12257 14565 12291
rect 14599 12288 14611 12291
rect 15286 12288 15292 12300
rect 14599 12260 15292 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12288 16083 12291
rect 16209 12291 16267 12297
rect 16209 12288 16221 12291
rect 16071 12260 16221 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 16209 12257 16221 12260
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 16945 12291 17003 12297
rect 16945 12288 16957 12291
rect 16724 12260 16957 12288
rect 16724 12248 16730 12260
rect 16945 12257 16957 12260
rect 16991 12288 17003 12291
rect 17218 12288 17224 12300
rect 16991 12260 17224 12288
rect 16991 12257 17003 12260
rect 16945 12251 17003 12257
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17635 12260 17969 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 13814 12180 13820 12232
rect 13872 12180 13878 12232
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 18046 12180 18052 12232
rect 18104 12180 18110 12232
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 14642 12152 14648 12164
rect 13740 12124 14648 12152
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 15286 12112 15292 12164
rect 15344 12112 15350 12164
rect 18524 12152 18552 12183
rect 17972 12124 18552 12152
rect 17972 12096 18000 12124
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12768 12056 12817 12084
rect 12768 12044 12774 12056
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 14182 12084 14188 12096
rect 13311 12056 14188 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 16850 12044 16856 12096
rect 16908 12044 16914 12096
rect 17954 12044 17960 12096
rect 18012 12044 18018 12096
rect 1104 11994 19228 12016
rect 1104 11942 3875 11994
rect 3927 11942 3939 11994
rect 3991 11942 4003 11994
rect 4055 11942 4067 11994
rect 4119 11942 4131 11994
rect 4183 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 8534 11994
rect 8586 11942 8598 11994
rect 8650 11942 8662 11994
rect 8714 11942 12937 11994
rect 12989 11942 13001 11994
rect 13053 11942 13065 11994
rect 13117 11942 13129 11994
rect 13181 11942 13193 11994
rect 13245 11942 17468 11994
rect 17520 11942 17532 11994
rect 17584 11942 17596 11994
rect 17648 11942 17660 11994
rect 17712 11942 17724 11994
rect 17776 11942 19228 11994
rect 1104 11920 19228 11942
rect 1670 11840 1676 11892
rect 1728 11840 1734 11892
rect 1946 11840 1952 11892
rect 2004 11840 2010 11892
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 1688 11812 1716 11840
rect 2148 11812 2176 11843
rect 4246 11840 4252 11892
rect 4304 11840 4310 11892
rect 6270 11840 6276 11892
rect 6328 11840 6334 11892
rect 8110 11840 8116 11892
rect 8168 11840 8174 11892
rect 8938 11840 8944 11892
rect 8996 11840 9002 11892
rect 9122 11840 9128 11892
rect 9180 11840 9186 11892
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 9858 11880 9864 11892
rect 9364 11852 9864 11880
rect 9364 11840 9370 11852
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 13078 11880 13084 11892
rect 11572 11852 13084 11880
rect 11572 11840 11578 11852
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 13725 11883 13783 11889
rect 13725 11849 13737 11883
rect 13771 11880 13783 11883
rect 13814 11880 13820 11892
rect 13771 11852 13820 11880
rect 13771 11849 13783 11852
rect 13725 11843 13783 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15344 11852 15393 11880
rect 15344 11840 15350 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 15381 11843 15439 11849
rect 15746 11840 15752 11892
rect 15804 11840 15810 11892
rect 16850 11840 16856 11892
rect 16908 11840 16914 11892
rect 2866 11812 2872 11824
rect 1688 11784 2176 11812
rect 2746 11784 2872 11812
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 2038 11744 2044 11756
rect 1903 11716 2044 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2314 11704 2320 11756
rect 2372 11704 2378 11756
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2746 11744 2774 11784
rect 2866 11772 2872 11784
rect 2924 11812 2930 11824
rect 3602 11812 3608 11824
rect 2924 11784 3608 11812
rect 2924 11772 2930 11784
rect 3602 11772 3608 11784
rect 3660 11772 3666 11824
rect 4982 11812 4988 11824
rect 3988 11784 4988 11812
rect 2455 11716 2774 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 3881 11747 3939 11753
rect 3881 11744 3893 11747
rect 3016 11716 3893 11744
rect 3016 11704 3022 11716
rect 3881 11713 3893 11716
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11645 2559 11679
rect 2501 11639 2559 11645
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 2639 11648 2789 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 2777 11645 2789 11648
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 2516 11540 2544 11639
rect 3050 11636 3056 11688
rect 3108 11676 3114 11688
rect 3988 11685 4016 11784
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6178 11744 6184 11756
rect 5859 11716 6184 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3108 11648 3341 11676
rect 3108 11636 3114 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4430 11676 4436 11688
rect 4304 11648 4436 11676
rect 4304 11636 4310 11648
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 4893 11679 4951 11685
rect 4893 11676 4905 11679
rect 4755 11648 4905 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 4893 11645 4905 11648
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5583 11648 5641 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11676 6055 11679
rect 6288 11676 6316 11840
rect 6914 11772 6920 11824
rect 6972 11812 6978 11824
rect 9140 11812 9168 11840
rect 6972 11784 7130 11812
rect 8312 11784 8800 11812
rect 6972 11772 6978 11784
rect 6362 11704 6368 11756
rect 6420 11704 6426 11756
rect 6043 11648 6316 11676
rect 6043 11645 6055 11648
rect 5997 11639 6055 11645
rect 2682 11568 2688 11620
rect 2740 11608 2746 11620
rect 3513 11611 3571 11617
rect 3513 11608 3525 11611
rect 2740 11580 3525 11608
rect 2740 11568 2746 11580
rect 3513 11577 3525 11580
rect 3559 11577 3571 11611
rect 3513 11571 3571 11577
rect 2774 11540 2780 11552
rect 2516 11512 2780 11540
rect 2774 11500 2780 11512
rect 2832 11540 2838 11552
rect 4632 11540 4660 11639
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 8312 11685 8340 11784
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 8435 11716 8708 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 2832 11512 4660 11540
rect 8680 11540 8708 11716
rect 8772 11676 8800 11784
rect 9140 11784 9628 11812
rect 9140 11744 9168 11784
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 9140 11716 9229 11744
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 9398 11704 9404 11756
rect 9456 11704 9462 11756
rect 9600 11753 9628 11784
rect 12158 11772 12164 11824
rect 12216 11812 12222 11824
rect 12253 11815 12311 11821
rect 12253 11812 12265 11815
rect 12216 11784 12265 11812
rect 12216 11772 12222 11784
rect 12253 11781 12265 11784
rect 12299 11781 12311 11815
rect 16298 11812 16304 11824
rect 12253 11775 12311 11781
rect 15580 11784 16304 11812
rect 15580 11756 15608 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9674 11704 9680 11756
rect 9732 11704 9738 11756
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 13354 11704 13360 11756
rect 13412 11704 13418 11756
rect 14182 11704 14188 11756
rect 14240 11704 14246 11756
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11744 15531 11747
rect 15562 11744 15568 11756
rect 15519 11716 15568 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16022 11744 16028 11756
rect 15979 11716 16028 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16868 11753 16896 11840
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16163 11716 16865 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8772 11648 9137 11676
rect 9125 11645 9137 11648
rect 9171 11676 9183 11679
rect 9692 11676 9720 11704
rect 9171 11648 9720 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11572 11648 11989 11676
rect 11572 11636 11578 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11676 14335 11679
rect 14642 11676 14648 11688
rect 14323 11648 14648 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 16040 11676 16068 11704
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 16040 11648 16773 11676
rect 16761 11645 16773 11648
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11608 8815 11611
rect 9398 11608 9404 11620
rect 8803 11580 9404 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 8680 11512 9689 11540
rect 2832 11500 2838 11512
rect 9677 11509 9689 11512
rect 9723 11509 9735 11543
rect 9677 11503 9735 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 12618 11540 12624 11552
rect 10836 11512 12624 11540
rect 10836 11500 10842 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 12952 11512 13829 11540
rect 12952 11500 12958 11512
rect 13817 11509 13829 11512
rect 13863 11509 13875 11543
rect 13817 11503 13875 11509
rect 1104 11450 19228 11472
rect 1104 11398 3215 11450
rect 3267 11398 3279 11450
rect 3331 11398 3343 11450
rect 3395 11398 3407 11450
rect 3459 11398 3471 11450
rect 3523 11398 7746 11450
rect 7798 11398 7810 11450
rect 7862 11398 7874 11450
rect 7926 11398 7938 11450
rect 7990 11398 8002 11450
rect 8054 11398 12277 11450
rect 12329 11398 12341 11450
rect 12393 11398 12405 11450
rect 12457 11398 12469 11450
rect 12521 11398 12533 11450
rect 12585 11398 16808 11450
rect 16860 11398 16872 11450
rect 16924 11398 16936 11450
rect 16988 11398 17000 11450
rect 17052 11398 17064 11450
rect 17116 11398 19228 11450
rect 1104 11376 19228 11398
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 3050 11336 3056 11348
rect 2639 11308 3056 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6638 11336 6644 11348
rect 6503 11308 6644 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 9766 11296 9772 11348
rect 9824 11296 9830 11348
rect 12158 11296 12164 11348
rect 12216 11296 12222 11348
rect 12894 11336 12900 11348
rect 12452 11308 12900 11336
rect 2958 11160 2964 11212
rect 3016 11160 3022 11212
rect 6638 11160 6644 11212
rect 6696 11160 6702 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6748 11172 7113 11200
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 4430 11132 4436 11144
rect 2823 11104 4436 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 6748 11141 6776 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7282 11200 7288 11212
rect 7101 11163 7159 11169
rect 7208 11172 7288 11200
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 7208 11141 7236 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7024 11064 7052 11092
rect 9784 11064 9812 11296
rect 11146 11268 11152 11280
rect 10704 11240 11152 11268
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 10594 11160 10600 11212
rect 10652 11160 10658 11212
rect 10704 11209 10732 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 12176 11268 12204 11296
rect 12253 11271 12311 11277
rect 12253 11268 12265 11271
rect 12176 11240 12265 11268
rect 12253 11237 12265 11240
rect 12299 11237 12311 11271
rect 12253 11231 12311 11237
rect 12452 11212 12480 11308
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 13412 11308 13461 11336
rect 13412 11296 13418 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 12710 11228 12716 11280
rect 12768 11228 12774 11280
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 11664 11172 12204 11200
rect 11664 11160 11670 11172
rect 9876 11132 9904 11160
rect 10778 11132 10784 11144
rect 9876 11104 10784 11132
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11146 11132 11152 11144
rect 10919 11104 11152 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12176 11132 12204 11172
rect 12434 11160 12440 11212
rect 12492 11160 12498 11212
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 12728 11141 12756 11228
rect 14918 11200 14924 11212
rect 13556 11172 14924 11200
rect 12529 11135 12587 11141
rect 12176 11104 12434 11132
rect 12069 11095 12127 11101
rect 7024 11036 9812 11064
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 12084 11064 12112 11095
rect 11112 11036 12112 11064
rect 12406 11064 12434 11104
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 12544 11064 12572 11095
rect 12912 11064 12940 11095
rect 13078 11092 13084 11144
rect 13136 11092 13142 11144
rect 13556 11141 13584 11172
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 12406 11036 12940 11064
rect 11112 11024 11118 11036
rect 10410 10956 10416 11008
rect 10468 10956 10474 11008
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 11517 10999 11575 11005
rect 11517 10996 11529 10999
rect 11296 10968 11529 10996
rect 11296 10956 11302 10968
rect 11517 10965 11529 10968
rect 11563 10965 11575 10999
rect 11517 10959 11575 10965
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 12989 10999 13047 11005
rect 12989 10996 13001 10999
rect 12768 10968 13001 10996
rect 12768 10956 12774 10968
rect 12989 10965 13001 10968
rect 13035 10965 13047 10999
rect 12989 10959 13047 10965
rect 18874 10956 18880 11008
rect 18932 10956 18938 11008
rect 1104 10906 19228 10928
rect 1104 10854 3875 10906
rect 3927 10854 3939 10906
rect 3991 10854 4003 10906
rect 4055 10854 4067 10906
rect 4119 10854 4131 10906
rect 4183 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 8534 10906
rect 8586 10854 8598 10906
rect 8650 10854 8662 10906
rect 8714 10854 12937 10906
rect 12989 10854 13001 10906
rect 13053 10854 13065 10906
rect 13117 10854 13129 10906
rect 13181 10854 13193 10906
rect 13245 10854 17468 10906
rect 17520 10854 17532 10906
rect 17584 10854 17596 10906
rect 17648 10854 17660 10906
rect 17712 10854 17724 10906
rect 17776 10854 19228 10906
rect 1104 10832 19228 10854
rect 4430 10752 4436 10804
rect 4488 10752 4494 10804
rect 10410 10792 10416 10804
rect 9600 10764 10416 10792
rect 9600 10733 9628 10764
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 11054 10752 11060 10804
rect 11112 10752 11118 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11204 10764 11529 10792
rect 11204 10752 11210 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 18322 10752 18328 10804
rect 18380 10792 18386 10804
rect 18417 10795 18475 10801
rect 18417 10792 18429 10795
rect 18380 10764 18429 10792
rect 18380 10752 18386 10764
rect 18417 10761 18429 10764
rect 18463 10761 18475 10795
rect 18417 10755 18475 10761
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10693 9643 10727
rect 11241 10727 11299 10733
rect 11241 10724 11253 10727
rect 10810 10696 11253 10724
rect 9585 10687 9643 10693
rect 11241 10693 11253 10696
rect 11287 10693 11299 10727
rect 15565 10727 15623 10733
rect 15565 10724 15577 10727
rect 11241 10687 11299 10693
rect 15212 10696 15577 10724
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 3988 10464 4016 10619
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 5169 10659 5227 10665
rect 5169 10656 5181 10659
rect 5092 10628 5181 10656
rect 5092 10600 5120 10628
rect 5169 10625 5181 10628
rect 5215 10656 5227 10659
rect 6454 10656 6460 10668
rect 5215 10628 6460 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 6454 10616 6460 10628
rect 6512 10656 6518 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6512 10628 6561 10656
rect 6512 10616 6518 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6822 10616 6828 10668
rect 6880 10616 6886 10668
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7524 10628 7757 10656
rect 7524 10616 7530 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11330 10665 11336 10668
rect 11325 10656 11336 10665
rect 11112 10628 11336 10656
rect 11112 10616 11118 10628
rect 11325 10619 11336 10628
rect 11330 10616 11336 10619
rect 11388 10616 11394 10668
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12710 10656 12716 10668
rect 12575 10628 12716 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 15212 10665 15240 10696
rect 15565 10693 15577 10696
rect 15611 10693 15623 10727
rect 15565 10687 15623 10693
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 16224 10656 16252 10752
rect 17678 10684 17684 10736
rect 17736 10684 17742 10736
rect 16482 10656 16488 10668
rect 15703 10628 16488 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4246 10588 4252 10600
rect 4111 10560 4252 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 5074 10548 5080 10600
rect 5132 10548 5138 10600
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7708 10560 7941 10588
rect 7708 10548 7714 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11296 10560 11897 10588
rect 11296 10548 11302 10560
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 12434 10548 12440 10600
rect 12492 10548 12498 10600
rect 15286 10548 15292 10600
rect 15344 10548 15350 10600
rect 16666 10548 16672 10600
rect 16724 10548 16730 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16776 10560 16957 10588
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10520 12955 10523
rect 13906 10520 13912 10532
rect 12943 10492 13912 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 16776 10520 16804 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 16632 10492 16804 10520
rect 16632 10480 16638 10492
rect 3970 10412 3976 10464
rect 4028 10412 4034 10464
rect 4246 10412 4252 10464
rect 4304 10412 4310 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 5224 10424 5273 10452
rect 5224 10412 5230 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 7558 10412 7564 10464
rect 7616 10412 7622 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14792 10424 14933 10452
rect 14792 10412 14798 10424
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 18509 10455 18567 10461
rect 18509 10452 18521 10455
rect 17552 10424 18521 10452
rect 17552 10412 17558 10424
rect 18509 10421 18521 10424
rect 18555 10421 18567 10455
rect 18509 10415 18567 10421
rect 1104 10362 19228 10384
rect 1104 10310 3215 10362
rect 3267 10310 3279 10362
rect 3331 10310 3343 10362
rect 3395 10310 3407 10362
rect 3459 10310 3471 10362
rect 3523 10310 7746 10362
rect 7798 10310 7810 10362
rect 7862 10310 7874 10362
rect 7926 10310 7938 10362
rect 7990 10310 8002 10362
rect 8054 10310 12277 10362
rect 12329 10310 12341 10362
rect 12393 10310 12405 10362
rect 12457 10310 12469 10362
rect 12521 10310 12533 10362
rect 12585 10310 16808 10362
rect 16860 10310 16872 10362
rect 16924 10310 16936 10362
rect 16988 10310 17000 10362
rect 17052 10310 17064 10362
rect 17116 10310 19228 10362
rect 1104 10288 19228 10310
rect 3970 10208 3976 10260
rect 4028 10208 4034 10260
rect 4246 10208 4252 10260
rect 4304 10208 4310 10260
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5040 10220 5917 10248
rect 5040 10208 5046 10220
rect 5905 10217 5917 10220
rect 5951 10217 5963 10251
rect 5905 10211 5963 10217
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 10505 10251 10563 10257
rect 7616 10220 7696 10248
rect 7616 10208 7622 10220
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 4154 10112 4160 10124
rect 3191 10084 4160 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 4264 10112 4292 10208
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4264 10084 4445 10112
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 6638 10072 6644 10124
rect 6696 10072 6702 10124
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7282 10112 7288 10124
rect 6779 10084 7288 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7668 10121 7696 10220
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10594 10248 10600 10260
rect 10551 10220 10600 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11756 10220 11989 10248
rect 11756 10208 11762 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15344 10220 16528 10248
rect 15344 10208 15350 10220
rect 16022 10140 16028 10192
rect 16080 10180 16086 10192
rect 16117 10183 16175 10189
rect 16117 10180 16129 10183
rect 16080 10152 16129 10180
rect 16080 10140 16086 10152
rect 16117 10149 16129 10152
rect 16163 10149 16175 10183
rect 16117 10143 16175 10149
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 11146 10112 11152 10124
rect 11011 10084 11152 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 14274 10072 14280 10124
rect 14332 10112 14338 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 14332 10084 14381 10112
rect 14332 10072 14338 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10112 14703 10115
rect 14734 10112 14740 10124
rect 14691 10084 14740 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 14734 10072 14740 10084
rect 14792 10072 14798 10124
rect 16500 10112 16528 10220
rect 16574 10208 16580 10260
rect 16632 10208 16638 10260
rect 17678 10208 17684 10260
rect 17736 10208 17742 10260
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 16500 10084 16773 10112
rect 16761 10081 16773 10084
rect 16807 10112 16819 10115
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 16807 10084 17877 10112
rect 16807 10081 16819 10084
rect 16761 10075 16819 10081
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10112 18199 10115
rect 18690 10112 18696 10124
rect 18187 10084 18696 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3421 10047 3479 10053
rect 3283 10016 3372 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 2130 9936 2136 9988
rect 2188 9936 2194 9988
rect 2866 9936 2872 9988
rect 2924 9936 2930 9988
rect 1394 9868 1400 9920
rect 1452 9868 1458 9920
rect 3234 9868 3240 9920
rect 3292 9868 3298 9920
rect 3344 9908 3372 10016
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3602 10044 3608 10056
rect 3467 10016 3608 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6963 10016 7113 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 3896 9908 3924 10007
rect 4080 9976 4108 10007
rect 4522 9976 4528 9988
rect 4080 9948 4528 9976
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 5166 9936 5172 9988
rect 5224 9936 5230 9988
rect 6840 9976 6868 10007
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8352 10016 8401 10044
rect 8352 10004 8358 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9030 10044 9036 10056
rect 8987 10016 9036 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 11238 10044 11244 10056
rect 10919 10016 11244 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10044 11483 10047
rect 11698 10044 11704 10056
rect 11471 10016 11704 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 13630 10044 13636 10056
rect 13311 10016 13636 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 16393 10047 16451 10053
rect 16393 10013 16405 10047
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 9214 9976 9220 9988
rect 6840 9948 9220 9976
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 11664 9948 12265 9976
rect 11664 9936 11670 9948
rect 12253 9945 12265 9948
rect 12299 9945 12311 9979
rect 16301 9979 16359 9985
rect 16301 9976 16313 9979
rect 15870 9948 16313 9976
rect 12253 9939 12311 9945
rect 16301 9945 16313 9948
rect 16347 9945 16359 9979
rect 16301 9939 16359 9945
rect 4798 9908 4804 9920
rect 3344 9880 4804 9908
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 6454 9868 6460 9920
rect 6512 9868 6518 9920
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7466 9908 7472 9920
rect 7064 9880 7472 9908
rect 7064 9868 7070 9880
rect 7466 9868 7472 9880
rect 7524 9908 7530 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7524 9880 7849 9908
rect 7524 9868 7530 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8996 9880 9045 9908
rect 8996 9868 9002 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 13814 9868 13820 9920
rect 13872 9868 13878 9920
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 16408 9908 16436 10007
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16540 10016 16865 10044
rect 16540 10004 16546 10016
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10044 17095 10047
rect 17494 10044 17500 10056
rect 17083 10016 17500 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 15620 9880 16436 9908
rect 15620 9868 15626 9880
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16960 9908 16988 10007
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 18322 10044 18328 10056
rect 18279 10016 18328 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 16540 9880 16988 9908
rect 17604 9908 17632 10007
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 17954 9908 17960 9920
rect 17604 9880 17960 9908
rect 16540 9868 16546 9880
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 1104 9818 19228 9840
rect 1104 9766 3875 9818
rect 3927 9766 3939 9818
rect 3991 9766 4003 9818
rect 4055 9766 4067 9818
rect 4119 9766 4131 9818
rect 4183 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 8534 9818
rect 8586 9766 8598 9818
rect 8650 9766 8662 9818
rect 8714 9766 12937 9818
rect 12989 9766 13001 9818
rect 13053 9766 13065 9818
rect 13117 9766 13129 9818
rect 13181 9766 13193 9818
rect 13245 9766 17468 9818
rect 17520 9766 17532 9818
rect 17584 9766 17596 9818
rect 17648 9766 17660 9818
rect 17712 9766 17724 9818
rect 17776 9766 19228 9818
rect 1104 9744 19228 9766
rect 2130 9664 2136 9716
rect 2188 9664 2194 9716
rect 2866 9664 2872 9716
rect 2924 9664 2930 9716
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 11204 9676 11529 9704
rect 11204 9664 11210 9676
rect 11517 9673 11529 9676
rect 11563 9673 11575 9707
rect 11517 9667 11575 9673
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 16482 9704 16488 9716
rect 15712 9676 16488 9704
rect 15712 9664 15718 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 18417 9707 18475 9713
rect 18417 9673 18429 9707
rect 18463 9704 18475 9707
rect 18690 9704 18696 9716
rect 18463 9676 18696 9704
rect 18463 9673 18475 9676
rect 18417 9667 18475 9673
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 5905 9639 5963 9645
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 5994 9636 6000 9648
rect 5951 9608 6000 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 8938 9596 8944 9648
rect 8996 9596 9002 9648
rect 9398 9596 9404 9648
rect 9456 9596 9462 9648
rect 11882 9636 11888 9648
rect 11348 9608 11888 9636
rect 2501 9571 2559 9577
rect 2041 9561 2099 9567
rect 2041 9527 2053 9561
rect 2087 9527 2099 9561
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 3234 9568 3240 9580
rect 2547 9540 3240 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4764 9540 4905 9568
rect 4764 9528 4770 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6822 9568 6828 9580
rect 6227 9540 6828 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 6963 9540 7205 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 7708 9540 7757 9568
rect 7708 9528 7714 9540
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11238 9568 11244 9580
rect 11195 9540 11244 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11348 9577 11376 9608
rect 11882 9596 11888 9608
rect 11940 9636 11946 9648
rect 14090 9636 14096 9648
rect 11940 9608 12434 9636
rect 13938 9608 14096 9636
rect 11940 9596 11946 9608
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 12406 9568 12434 9608
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14274 9596 14280 9648
rect 14332 9636 14338 9648
rect 18601 9639 18659 9645
rect 18601 9636 18613 9639
rect 14332 9608 15424 9636
rect 18170 9608 18613 9636
rect 14332 9596 14338 9608
rect 14660 9580 14688 9608
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12406 9540 12541 9568
rect 11333 9531 11391 9537
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 14642 9528 14648 9580
rect 14700 9528 14706 9580
rect 14734 9528 14740 9580
rect 14792 9528 14798 9580
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14976 9540 15025 9568
rect 14976 9528 14982 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15396 9568 15424 9608
rect 18601 9605 18613 9608
rect 18647 9605 18659 9639
rect 18601 9599 18659 9605
rect 16666 9568 16672 9580
rect 15396 9540 16672 9568
rect 15013 9531 15071 9537
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 2041 9521 2099 9527
rect 2056 9444 2084 9521
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2372 9472 2421 9500
rect 2372 9460 2378 9472
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9500 6607 9503
rect 6638 9500 6644 9512
rect 6595 9472 6644 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 2038 9392 2044 9444
rect 2096 9432 2102 9444
rect 5092 9432 5120 9460
rect 2096 9404 5120 9432
rect 2096 9392 2102 9404
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5074 9364 5080 9376
rect 4856 9336 5080 9364
rect 4856 9324 4862 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 6840 9364 6868 9528
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 11514 9500 11520 9512
rect 9723 9472 11520 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 12161 9503 12219 9509
rect 12161 9500 12173 9503
rect 11756 9472 12173 9500
rect 11756 9460 11762 9472
rect 12161 9469 12173 9472
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12483 9472 12517 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9432 7987 9435
rect 8294 9432 8300 9444
rect 7975 9404 8300 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 11146 9392 11152 9444
rect 11204 9432 11210 9444
rect 12452 9432 12480 9463
rect 12710 9460 12716 9512
rect 12768 9460 12774 9512
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 13964 9472 14381 9500
rect 13964 9460 13970 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 16206 9460 16212 9512
rect 16264 9500 16270 9512
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16264 9472 16957 9500
rect 16264 9460 16270 9472
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18524 9500 18552 9531
rect 18012 9472 18552 9500
rect 18012 9460 18018 9472
rect 13354 9432 13360 9444
rect 11204 9404 13360 9432
rect 11204 9392 11210 9404
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 9214 9364 9220 9376
rect 6840 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 11238 9324 11244 9376
rect 11296 9324 11302 9376
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12253 9367 12311 9373
rect 12253 9364 12265 9367
rect 12032 9336 12265 9364
rect 12032 9324 12038 9336
rect 12253 9333 12265 9336
rect 12299 9333 12311 9367
rect 12253 9327 12311 9333
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13630 9364 13636 9376
rect 12943 9336 13636 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 1104 9274 19228 9296
rect 1104 9222 3215 9274
rect 3267 9222 3279 9274
rect 3331 9222 3343 9274
rect 3395 9222 3407 9274
rect 3459 9222 3471 9274
rect 3523 9222 7746 9274
rect 7798 9222 7810 9274
rect 7862 9222 7874 9274
rect 7926 9222 7938 9274
rect 7990 9222 8002 9274
rect 8054 9222 12277 9274
rect 12329 9222 12341 9274
rect 12393 9222 12405 9274
rect 12457 9222 12469 9274
rect 12521 9222 12533 9274
rect 12585 9222 16808 9274
rect 16860 9222 16872 9274
rect 16924 9222 16936 9274
rect 16988 9222 17000 9274
rect 17052 9222 17064 9274
rect 17116 9222 19228 9274
rect 1104 9200 19228 9222
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7708 9132 8033 9160
rect 7708 9120 7714 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 8021 9123 8079 9129
rect 11146 9120 11152 9172
rect 11204 9120 11210 9172
rect 11238 9120 11244 9172
rect 11296 9120 11302 9172
rect 12621 9163 12679 9169
rect 12621 9129 12633 9163
rect 12667 9160 12679 9163
rect 12710 9160 12716 9172
rect 12667 9132 12716 9160
rect 12667 9129 12679 9132
rect 12621 9123 12679 9129
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 13354 9120 13360 9172
rect 13412 9120 13418 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 14148 9132 14657 9160
rect 14148 9120 14154 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 16117 9163 16175 9169
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16206 9160 16212 9172
rect 16163 9132 16212 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1452 8996 1961 9024
rect 1452 8984 1458 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2406 8984 2412 9036
rect 2464 8984 2470 9036
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 9024 6331 9027
rect 6638 9024 6644 9036
rect 6319 8996 6644 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 11164 9033 11192 9120
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1964 8928 2053 8956
rect 1964 8832 1992 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2498 8916 2504 8968
rect 2556 8916 2562 8968
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 4982 8956 4988 8968
rect 2832 8928 4988 8956
rect 2832 8916 2838 8928
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8956 9091 8959
rect 9214 8956 9220 8968
rect 9079 8928 9220 8956
rect 9079 8925 9091 8928
rect 9033 8919 9091 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8956 9367 8959
rect 9398 8956 9404 8968
rect 9355 8928 9404 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 9398 8916 9404 8928
rect 9456 8956 9462 8968
rect 10962 8956 10968 8968
rect 9456 8928 10968 8956
rect 9456 8916 9462 8928
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11256 8956 11284 9120
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 14461 9027 14519 9033
rect 14461 9024 14473 9027
rect 13740 8996 14473 9024
rect 11103 8928 11284 8956
rect 13265 8959 13323 8965
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 13265 8925 13277 8959
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 6454 8848 6460 8900
rect 6512 8888 6518 8900
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 6512 8860 6561 8888
rect 6512 8848 6518 8860
rect 6549 8857 6561 8860
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 7006 8848 7012 8900
rect 7064 8848 7070 8900
rect 13280 8888 13308 8919
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13740 8965 13768 8996
rect 14461 8993 14473 8996
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16574 9024 16580 9036
rect 15979 8996 16580 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13596 8928 13737 8956
rect 13596 8916 13602 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13872 8928 14289 8956
rect 13872 8916 13878 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 14918 8956 14924 8968
rect 14783 8928 14924 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 15838 8916 15844 8968
rect 15896 8916 15902 8968
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 17862 8956 17868 8968
rect 16448 8928 17868 8956
rect 16448 8916 16454 8928
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 14093 8891 14151 8897
rect 14093 8888 14105 8891
rect 13280 8860 14105 8888
rect 14093 8857 14105 8860
rect 14139 8857 14151 8891
rect 14093 8851 14151 8857
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 3016 8792 3157 8820
rect 3016 8780 3022 8792
rect 3145 8789 3157 8792
rect 3191 8789 3203 8823
rect 3145 8783 3203 8789
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 10134 8820 10140 8832
rect 4764 8792 10140 8820
rect 4764 8780 4770 8792
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 10686 8780 10692 8832
rect 10744 8780 10750 8832
rect 1104 8730 19228 8752
rect 1104 8678 3875 8730
rect 3927 8678 3939 8730
rect 3991 8678 4003 8730
rect 4055 8678 4067 8730
rect 4119 8678 4131 8730
rect 4183 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 8534 8730
rect 8586 8678 8598 8730
rect 8650 8678 8662 8730
rect 8714 8678 12937 8730
rect 12989 8678 13001 8730
rect 13053 8678 13065 8730
rect 13117 8678 13129 8730
rect 13181 8678 13193 8730
rect 13245 8678 17468 8730
rect 17520 8678 17532 8730
rect 17584 8678 17596 8730
rect 17648 8678 17660 8730
rect 17712 8678 17724 8730
rect 17776 8678 19228 8730
rect 1104 8656 19228 8678
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 5166 8616 5172 8628
rect 4172 8588 5172 8616
rect 2424 8480 2452 8576
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 3528 8520 4077 8548
rect 3528 8489 3556 8520
rect 4065 8517 4077 8520
rect 4111 8517 4123 8551
rect 4065 8511 4123 8517
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2424 8452 2697 8480
rect 2685 8449 2697 8452
rect 2731 8480 2743 8483
rect 2976 8480 3096 8486
rect 2731 8458 3096 8480
rect 2731 8452 3004 8458
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 2004 8384 2329 8412
rect 2004 8372 2010 8384
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 2792 8344 2820 8375
rect 2866 8372 2872 8424
rect 2924 8372 2930 8424
rect 2958 8372 2964 8424
rect 3016 8372 3022 8424
rect 3068 8412 3096 8458
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4172 8489 4200 8588
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 7006 8576 7012 8628
rect 7064 8576 7070 8628
rect 10686 8616 10692 8628
rect 9416 8588 10692 8616
rect 5534 8508 5540 8560
rect 5592 8508 5598 8560
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3844 8452 3985 8480
rect 3844 8440 3850 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 6012 8480 6040 8576
rect 9306 8548 9312 8560
rect 9140 8520 9312 8548
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6012 8452 6929 8480
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 9140 8489 9168 8520
rect 9306 8508 9312 8520
rect 9364 8508 9370 8560
rect 9416 8557 9444 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10873 8619 10931 8625
rect 10873 8585 10885 8619
rect 10919 8616 10931 8619
rect 11698 8616 11704 8628
rect 10919 8588 11704 8616
rect 10919 8585 10931 8588
rect 10873 8579 10931 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11974 8616 11980 8628
rect 11808 8588 11980 8616
rect 9401 8551 9459 8557
rect 9401 8517 9413 8551
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 9858 8508 9864 8560
rect 9916 8508 9922 8560
rect 11808 8557 11836 8588
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 13538 8616 13544 8628
rect 13311 8588 13544 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14642 8576 14648 8628
rect 14700 8576 14706 8628
rect 18506 8616 18512 8628
rect 16040 8588 18512 8616
rect 11793 8551 11851 8557
rect 11793 8517 11805 8551
rect 11839 8517 11851 8551
rect 11793 8511 11851 8517
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 8352 8452 9137 8480
rect 8352 8440 8358 8452
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 12894 8440 12900 8492
rect 12952 8440 12958 8492
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8449 13415 8483
rect 13357 8443 13415 8449
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3068 8384 3433 8412
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 3804 8344 3832 8440
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 3896 8384 4537 8412
rect 3896 8353 3924 8384
rect 4525 8381 4537 8384
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 11514 8372 11520 8424
rect 11572 8372 11578 8424
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 13372 8412 13400 8443
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 14734 8480 14740 8492
rect 13872 8452 14740 8480
rect 13872 8440 13878 8452
rect 14734 8440 14740 8452
rect 14792 8480 14798 8492
rect 16040 8489 16068 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 16482 8548 16488 8560
rect 16132 8520 16488 8548
rect 15197 8483 15255 8489
rect 15197 8480 15209 8483
rect 14792 8452 15209 8480
rect 14792 8440 14798 8452
rect 15197 8449 15209 8452
rect 15243 8449 15255 8483
rect 15197 8443 15255 8449
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 12860 8384 13400 8412
rect 12860 8372 12866 8384
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15562 8412 15568 8424
rect 15519 8384 15568 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15562 8372 15568 8384
rect 15620 8372 15626 8424
rect 16132 8421 16160 8520
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 17402 8508 17408 8560
rect 17460 8508 17466 8560
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8480 16267 8483
rect 16390 8480 16396 8492
rect 16255 8452 16396 8480
rect 16255 8449 16267 8452
rect 16209 8443 16267 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8381 16175 8415
rect 16117 8375 16175 8381
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 16945 8415 17003 8421
rect 16945 8412 16957 8415
rect 16531 8384 16957 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 16945 8381 16957 8384
rect 16991 8381 17003 8415
rect 16945 8375 17003 8381
rect 2547 8316 2728 8344
rect 2792 8316 3832 8344
rect 3881 8347 3939 8353
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 1762 8236 1768 8288
rect 1820 8236 1826 8288
rect 2700 8276 2728 8316
rect 3881 8313 3893 8347
rect 3927 8313 3939 8347
rect 15304 8344 15332 8372
rect 16132 8344 16160 8375
rect 3881 8307 3939 8313
rect 5920 8316 6132 8344
rect 15304 8316 16160 8344
rect 16316 8344 16344 8375
rect 16574 8344 16580 8356
rect 16316 8316 16580 8344
rect 2866 8276 2872 8288
rect 2700 8248 2872 8276
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5920 8276 5948 8316
rect 5132 8248 5948 8276
rect 5132 8236 5138 8248
rect 5994 8236 6000 8288
rect 6052 8236 6058 8288
rect 6104 8276 6132 8316
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 8754 8276 8760 8288
rect 6104 8248 8760 8276
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 16592 8276 16620 8304
rect 17586 8276 17592 8288
rect 16592 8248 17592 8276
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 18414 8236 18420 8288
rect 18472 8236 18478 8288
rect 1104 8186 19228 8208
rect 1104 8134 3215 8186
rect 3267 8134 3279 8186
rect 3331 8134 3343 8186
rect 3395 8134 3407 8186
rect 3459 8134 3471 8186
rect 3523 8134 7746 8186
rect 7798 8134 7810 8186
rect 7862 8134 7874 8186
rect 7926 8134 7938 8186
rect 7990 8134 8002 8186
rect 8054 8134 12277 8186
rect 12329 8134 12341 8186
rect 12393 8134 12405 8186
rect 12457 8134 12469 8186
rect 12521 8134 12533 8186
rect 12585 8134 16808 8186
rect 16860 8134 16872 8186
rect 16924 8134 16936 8186
rect 16988 8134 17000 8186
rect 17052 8134 17064 8186
rect 17116 8134 19228 8186
rect 1104 8112 19228 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 2498 8072 2504 8084
rect 1811 8044 2504 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 4338 8032 4344 8084
rect 4396 8032 4402 8084
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 5534 8072 5540 8084
rect 4479 8044 5540 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 9493 8075 9551 8081
rect 7576 8044 8524 8072
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1762 7936 1768 7948
rect 1443 7908 1768 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 4356 7936 4384 8032
rect 7576 8004 7604 8044
rect 4724 7976 7604 8004
rect 4724 7936 4752 7976
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 7708 7976 7849 8004
rect 7708 7964 7714 7976
rect 7837 7973 7849 7976
rect 7883 7973 7895 8007
rect 7837 7967 7895 7973
rect 4356 7908 4752 7936
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1412 7840 1593 7868
rect 1412 7812 1440 7840
rect 1581 7837 1593 7840
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 4154 7868 4160 7880
rect 3651 7840 4160 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 4724 7868 4752 7908
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 7926 7936 7932 7948
rect 4847 7908 7932 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 7926 7896 7932 7908
rect 7984 7936 7990 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7984 7908 8125 7936
rect 7984 7896 7990 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4724 7840 4905 7868
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 8496 7877 8524 8044
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9858 8072 9864 8084
rect 9539 8044 9864 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11514 8072 11520 8084
rect 10919 8044 11520 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 12802 8072 12808 8084
rect 12176 8044 12808 8072
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 8812 7908 11652 7936
rect 8812 7896 8818 7908
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8481 7871 8539 7877
rect 8251 7840 8432 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 1394 7760 1400 7812
rect 1452 7760 1458 7812
rect 4172 7800 4200 7828
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 4172 7772 5273 7800
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 5261 7763 5319 7769
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 7006 7800 7012 7812
rect 6696 7772 7012 7800
rect 6696 7760 6702 7772
rect 7006 7760 7012 7772
rect 7064 7800 7070 7812
rect 8404 7800 8432 7840
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8772 7868 8800 7896
rect 11624 7880 11652 7908
rect 8711 7840 8800 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 9398 7828 9404 7880
rect 9456 7828 9462 7880
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11606 7828 11612 7880
rect 11664 7828 11670 7880
rect 12176 7877 12204 8044
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 15378 8072 15384 8084
rect 15028 8044 15384 8072
rect 12345 8007 12403 8013
rect 12345 7973 12357 8007
rect 12391 8004 12403 8007
rect 12894 8004 12900 8016
rect 12391 7976 12900 8004
rect 12391 7973 12403 7976
rect 12345 7967 12403 7973
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 13587 7908 14749 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 14737 7905 14749 7908
rect 14783 7936 14795 7939
rect 14918 7936 14924 7948
rect 14783 7908 14924 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 15028 7945 15056 8044
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 17310 8032 17316 8084
rect 17368 8032 17374 8084
rect 17402 8032 17408 8084
rect 17460 8032 17466 8084
rect 17586 8032 17592 8084
rect 17644 8032 17650 8084
rect 15120 7976 15700 8004
rect 15013 7939 15071 7945
rect 15013 7905 15025 7939
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 13998 7868 14004 7880
rect 13771 7840 14004 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 8573 7803 8631 7809
rect 8573 7800 8585 7803
rect 7064 7772 8248 7800
rect 8404 7772 8585 7800
rect 7064 7760 7070 7772
rect 8220 7744 8248 7772
rect 8573 7769 8585 7772
rect 8619 7769 8631 7803
rect 11072 7800 11100 7828
rect 12268 7800 12296 7831
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 15120 7877 15148 7976
rect 15672 7936 15700 7976
rect 17328 7936 17356 8032
rect 18064 7976 18828 8004
rect 18064 7945 18092 7976
rect 18800 7948 18828 7976
rect 15672 7908 17356 7936
rect 18049 7939 18107 7945
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15194 7828 15200 7880
rect 15252 7828 15258 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15470 7868 15476 7880
rect 15289 7831 15347 7837
rect 15396 7840 15476 7868
rect 11072 7772 12296 7800
rect 13909 7803 13967 7809
rect 8573 7763 8631 7769
rect 13909 7769 13921 7803
rect 13955 7800 13967 7803
rect 15304 7800 15332 7831
rect 13955 7772 15332 7800
rect 15396 7800 15424 7840
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15672 7877 15700 7908
rect 18049 7905 18061 7939
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7936 18383 7939
rect 18414 7936 18420 7948
rect 18371 7908 18420 7936
rect 18371 7905 18383 7908
rect 18325 7899 18383 7905
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7868 15991 7871
rect 16390 7868 16396 7880
rect 15979 7840 16396 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 15764 7800 15792 7831
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7837 17371 7871
rect 17313 7831 17371 7837
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7868 18015 7871
rect 18340 7868 18368 7899
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 18782 7896 18788 7948
rect 18840 7896 18846 7948
rect 18003 7840 18368 7868
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 15396 7772 15792 7800
rect 17328 7800 17356 7831
rect 17862 7800 17868 7812
rect 17328 7772 17868 7800
rect 13955 7769 13967 7772
rect 13909 7763 13967 7769
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 3142 7732 3148 7744
rect 2372 7704 3148 7732
rect 2372 7692 2378 7704
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 4614 7692 4620 7744
rect 4672 7692 4678 7744
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 8202 7692 8208 7744
rect 8260 7692 8266 7744
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 10410 7732 10416 7744
rect 10192 7704 10416 7732
rect 10192 7692 10198 7704
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 14826 7692 14832 7744
rect 14884 7692 14890 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15396 7732 15424 7772
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 15252 7704 15424 7732
rect 15252 7692 15258 7704
rect 15470 7692 15476 7744
rect 15528 7692 15534 7744
rect 18877 7735 18935 7741
rect 18877 7701 18889 7735
rect 18923 7732 18935 7735
rect 18923 7704 19288 7732
rect 18923 7701 18935 7704
rect 18877 7695 18935 7701
rect 1104 7642 19228 7664
rect 1104 7590 3875 7642
rect 3927 7590 3939 7642
rect 3991 7590 4003 7642
rect 4055 7590 4067 7642
rect 4119 7590 4131 7642
rect 4183 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 8534 7642
rect 8586 7590 8598 7642
rect 8650 7590 8662 7642
rect 8714 7590 12937 7642
rect 12989 7590 13001 7642
rect 13053 7590 13065 7642
rect 13117 7590 13129 7642
rect 13181 7590 13193 7642
rect 13245 7590 17468 7642
rect 17520 7590 17532 7642
rect 17584 7590 17596 7642
rect 17648 7590 17660 7642
rect 17712 7590 17724 7642
rect 17776 7590 19228 7642
rect 1104 7568 19228 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 1946 7528 1952 7540
rect 1443 7500 1952 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 4614 7528 4620 7540
rect 4448 7500 4620 7528
rect 2222 7420 2228 7472
rect 2280 7420 2286 7472
rect 2866 7420 2872 7472
rect 2924 7420 2930 7472
rect 4264 7460 4292 7488
rect 4448 7469 4476 7500
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 5132 7500 7021 7528
rect 5132 7488 5138 7500
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 7009 7491 7067 7497
rect 7098 7488 7104 7540
rect 7156 7488 7162 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 9674 7488 9680 7540
rect 9732 7488 9738 7540
rect 10134 7488 10140 7540
rect 10192 7488 10198 7540
rect 10410 7488 10416 7540
rect 10468 7488 10474 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 14090 7528 14096 7540
rect 13679 7500 14096 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 14826 7488 14832 7540
rect 14884 7488 14890 7540
rect 14918 7488 14924 7540
rect 14976 7488 14982 7540
rect 17126 7488 17132 7540
rect 17184 7488 17190 7540
rect 18506 7488 18512 7540
rect 18564 7488 18570 7540
rect 4172 7432 4292 7460
rect 4433 7463 4491 7469
rect 3142 7352 3148 7404
rect 3200 7392 3206 7404
rect 4172 7401 4200 7432
rect 4433 7429 4445 7463
rect 4479 7429 4491 7463
rect 4433 7423 4491 7429
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3200 7364 4169 7392
rect 3200 7352 3206 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 5920 7364 6745 7392
rect 5920 7333 5948 7364
rect 6733 7361 6745 7364
rect 6779 7392 6791 7395
rect 7116 7392 7144 7488
rect 6779 7364 7144 7392
rect 7193 7395 7251 7401
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7760 7392 7788 7488
rect 8220 7460 8248 7488
rect 7944 7432 8248 7460
rect 7944 7401 7972 7432
rect 8938 7420 8944 7472
rect 8996 7420 9002 7472
rect 7423 7364 7788 7392
rect 7929 7395 7987 7401
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 9692 7392 9720 7488
rect 10318 7460 10324 7472
rect 10060 7432 10324 7460
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9692 7364 9965 7392
rect 7929 7355 7987 7361
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6052 7296 6653 7324
rect 6052 7284 6058 7296
rect 6641 7293 6653 7296
rect 6687 7324 6699 7327
rect 7208 7324 7236 7355
rect 6687 7296 7236 7324
rect 8205 7327 8263 7333
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 9398 7324 9404 7336
rect 8251 7296 9404 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 9398 7284 9404 7296
rect 9456 7324 9462 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9456 7296 9781 7324
rect 9456 7284 9462 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 7926 7216 7932 7268
rect 7984 7216 7990 7268
rect 9677 7259 9735 7265
rect 9677 7225 9689 7259
rect 9723 7256 9735 7259
rect 10060 7256 10088 7432
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 10428 7460 10456 7488
rect 10428 7432 10640 7460
rect 10612 7404 10640 7432
rect 12894 7420 12900 7472
rect 12952 7420 12958 7472
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10275 7390 10364 7392
rect 10428 7390 10517 7392
rect 10275 7364 10517 7390
rect 10275 7361 10287 7364
rect 10336 7362 10456 7364
rect 10229 7355 10287 7361
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 10520 7324 10548 7355
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11514 7392 11520 7404
rect 11020 7364 11520 7392
rect 11020 7352 11026 7364
rect 11514 7352 11520 7364
rect 11572 7392 11578 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11572 7364 11897 7392
rect 11572 7352 11578 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 14844 7392 14872 7488
rect 14936 7401 14964 7488
rect 11885 7355 11943 7361
rect 13648 7364 14872 7392
rect 14921 7395 14979 7401
rect 12161 7327 12219 7333
rect 10520 7296 10640 7324
rect 9723 7228 10088 7256
rect 9723 7225 9735 7228
rect 9677 7219 9735 7225
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7188 6423 7191
rect 7944 7188 7972 7216
rect 6411 7160 7972 7188
rect 6411 7157 6423 7160
rect 6365 7151 6423 7157
rect 10410 7148 10416 7200
rect 10468 7148 10474 7200
rect 10612 7188 10640 7296
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 13648 7324 13676 7364
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 15252 7364 16681 7392
rect 15252 7352 15258 7364
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 17144 7392 17172 7488
rect 16899 7364 17172 7392
rect 18693 7395 18751 7401
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 18782 7392 18788 7404
rect 18739 7364 18788 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 12207 7296 13676 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 14090 7284 14096 7336
rect 14148 7284 14154 7336
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7324 14703 7327
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14691 7296 14841 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 15378 7324 15384 7336
rect 15335 7296 15384 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16868 7324 16896 7355
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19260 7392 19288 7704
rect 18923 7364 19288 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 16632 7296 16896 7324
rect 16632 7284 16638 7296
rect 15580 7228 18644 7256
rect 15580 7188 15608 7228
rect 18616 7200 18644 7228
rect 10612 7160 15608 7188
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 16724 7160 16773 7188
rect 16724 7148 16730 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 18598 7148 18604 7200
rect 18656 7148 18662 7200
rect 1104 7098 19228 7120
rect 1104 7046 3215 7098
rect 3267 7046 3279 7098
rect 3331 7046 3343 7098
rect 3395 7046 3407 7098
rect 3459 7046 3471 7098
rect 3523 7046 7746 7098
rect 7798 7046 7810 7098
rect 7862 7046 7874 7098
rect 7926 7046 7938 7098
rect 7990 7046 8002 7098
rect 8054 7046 12277 7098
rect 12329 7046 12341 7098
rect 12393 7046 12405 7098
rect 12457 7046 12469 7098
rect 12521 7046 12533 7098
rect 12585 7046 16808 7098
rect 16860 7046 16872 7098
rect 16924 7046 16936 7098
rect 16988 7046 17000 7098
rect 17052 7046 17064 7098
rect 17116 7046 19228 7098
rect 1104 7024 19228 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2317 6987 2375 6993
rect 2317 6984 2329 6987
rect 2280 6956 2329 6984
rect 2280 6944 2286 6956
rect 2317 6953 2329 6956
rect 2363 6953 2375 6987
rect 2317 6947 2375 6953
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4246 6984 4252 6996
rect 4203 6956 4252 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4246 6944 4252 6956
rect 4304 6984 4310 6996
rect 4982 6984 4988 6996
rect 4304 6956 4988 6984
rect 4304 6944 4310 6956
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 8938 6944 8944 6996
rect 8996 6984 9002 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8996 6956 9045 6984
rect 8996 6944 9002 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 9033 6947 9091 6953
rect 10594 6944 10600 6996
rect 10652 6944 10658 6996
rect 12894 6944 12900 6996
rect 12952 6944 12958 6996
rect 13998 6944 14004 6996
rect 14056 6984 14062 6996
rect 14185 6987 14243 6993
rect 14185 6984 14197 6987
rect 14056 6956 14197 6984
rect 14056 6944 14062 6956
rect 14185 6953 14197 6956
rect 14231 6953 14243 6987
rect 14185 6947 14243 6953
rect 10612 6916 10640 6944
rect 15194 6916 15200 6928
rect 10612 6888 15200 6916
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2590 6848 2596 6860
rect 1912 6820 2596 6848
rect 1912 6808 1918 6820
rect 2590 6808 2596 6820
rect 2648 6848 2654 6860
rect 5166 6848 5172 6860
rect 2648 6820 2774 6848
rect 2648 6808 2654 6820
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2746 6780 2774 6820
rect 4908 6820 5172 6848
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2746 6752 2973 6780
rect 2225 6743 2283 6749
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3191 6752 3924 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 2240 6712 2268 6743
rect 2682 6712 2688 6724
rect 2240 6684 2688 6712
rect 2682 6672 2688 6684
rect 2740 6712 2746 6724
rect 3896 6721 3924 6752
rect 3881 6715 3939 6721
rect 2740 6684 3832 6712
rect 2740 6672 2746 6684
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 3804 6644 3832 6684
rect 3881 6681 3893 6715
rect 3927 6712 3939 6715
rect 4908 6712 4936 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9398 6848 9404 6860
rect 9355 6820 9404 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5534 6780 5540 6792
rect 5123 6752 5540 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 3927 6684 4936 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 4338 6644 4344 6656
rect 3804 6616 4344 6644
rect 4338 6604 4344 6616
rect 4396 6644 4402 6656
rect 5000 6644 5028 6743
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8772 6752 8953 6780
rect 8772 6656 8800 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 10410 6780 10416 6792
rect 9539 6752 10416 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11606 6740 11612 6792
rect 11664 6740 11670 6792
rect 12268 6789 12296 6888
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 15286 6876 15292 6928
rect 15344 6916 15350 6928
rect 15344 6888 16252 6916
rect 15344 6876 15350 6888
rect 13722 6848 13728 6860
rect 12820 6820 13728 6848
rect 12820 6792 12848 6820
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 15304 6848 15332 6876
rect 15212 6820 15332 6848
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11808 6752 12081 6780
rect 11808 6656 11836 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14148 6752 14749 6780
rect 14148 6740 14154 6752
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 11977 6715 12035 6721
rect 11977 6681 11989 6715
rect 12023 6712 12035 6715
rect 15212 6712 15240 6820
rect 15378 6808 15384 6860
rect 15436 6808 15442 6860
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 15470 6780 15476 6792
rect 15335 6752 15476 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 16025 6783 16083 6789
rect 15620 6752 15976 6780
rect 15620 6740 15626 6752
rect 15948 6724 15976 6752
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 12023 6684 15240 6712
rect 12023 6681 12035 6684
rect 11977 6675 12035 6681
rect 15930 6672 15936 6724
rect 15988 6672 15994 6724
rect 16040 6656 16068 6743
rect 5442 6644 5448 6656
rect 4396 6616 5448 6644
rect 4396 6604 4402 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 8754 6604 8760 6656
rect 8812 6604 8818 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 11790 6604 11796 6656
rect 11848 6604 11854 6656
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6644 12311 6647
rect 12618 6644 12624 6656
rect 12299 6616 12624 6644
rect 12299 6613 12311 6616
rect 12253 6607 12311 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 14918 6604 14924 6656
rect 14976 6604 14982 6656
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15657 6647 15715 6653
rect 15657 6644 15669 6647
rect 15620 6616 15669 6644
rect 15620 6604 15626 6616
rect 15657 6613 15669 6616
rect 15703 6613 15715 6647
rect 15657 6607 15715 6613
rect 15838 6604 15844 6656
rect 15896 6604 15902 6656
rect 16022 6604 16028 6656
rect 16080 6604 16086 6656
rect 16132 6644 16160 6811
rect 16224 6789 16252 6888
rect 16850 6808 16856 6860
rect 16908 6848 16914 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 16908 6820 17877 6848
rect 16908 6808 16914 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 16347 6752 16589 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 16758 6740 16764 6792
rect 16816 6780 16822 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 16816 6752 17141 6780
rect 16816 6740 16822 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 16574 6644 16580 6656
rect 16132 6616 16580 6644
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 17313 6647 17371 6653
rect 17313 6644 17325 6647
rect 17092 6616 17325 6644
rect 17092 6604 17098 6616
rect 17313 6613 17325 6616
rect 17359 6613 17371 6647
rect 17313 6607 17371 6613
rect 1104 6554 19228 6576
rect 1104 6502 3875 6554
rect 3927 6502 3939 6554
rect 3991 6502 4003 6554
rect 4055 6502 4067 6554
rect 4119 6502 4131 6554
rect 4183 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 8534 6554
rect 8586 6502 8598 6554
rect 8650 6502 8662 6554
rect 8714 6502 12937 6554
rect 12989 6502 13001 6554
rect 13053 6502 13065 6554
rect 13117 6502 13129 6554
rect 13181 6502 13193 6554
rect 13245 6502 17468 6554
rect 17520 6502 17532 6554
rect 17584 6502 17596 6554
rect 17648 6502 17660 6554
rect 17712 6502 17724 6554
rect 17776 6502 19228 6554
rect 1104 6480 19228 6502
rect 3050 6400 3056 6452
rect 3108 6400 3114 6452
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 3200 6412 3648 6440
rect 3200 6400 3206 6412
rect 2222 6332 2228 6384
rect 2280 6332 2286 6384
rect 3068 6372 3096 6400
rect 3068 6344 3188 6372
rect 3160 6313 3188 6344
rect 3620 6313 3648 6412
rect 5166 6400 5172 6452
rect 5224 6400 5230 6452
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 14700 6412 17172 6440
rect 14700 6400 14706 6412
rect 5184 6372 5212 6400
rect 4632 6344 5212 6372
rect 7377 6375 7435 6381
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6304 4583 6307
rect 4632 6304 4660 6344
rect 7377 6341 7389 6375
rect 7423 6372 7435 6375
rect 7650 6372 7656 6384
rect 7423 6344 7656 6372
rect 7423 6341 7435 6344
rect 7377 6335 7435 6341
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 9490 6372 9496 6384
rect 8602 6344 9496 6372
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 4571 6276 4660 6304
rect 4709 6307 4767 6313
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6236 2927 6239
rect 3697 6239 3755 6245
rect 2915 6208 3280 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 3252 6177 3280 6208
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 3786 6236 3792 6248
rect 3743 6208 3792 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 4724 6236 4752 6267
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 7064 6276 7113 6304
rect 7064 6264 7070 6276
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 9692 6304 9720 6400
rect 12802 6372 12808 6384
rect 10612 6344 12808 6372
rect 10612 6313 10640 6344
rect 12802 6332 12808 6344
rect 12860 6332 12866 6384
rect 14660 6372 14688 6400
rect 14568 6344 14688 6372
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9692 6276 9873 6304
rect 7101 6267 7159 6273
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 5258 6236 5264 6248
rect 4540 6208 5264 6236
rect 3237 6171 3295 6177
rect 3237 6137 3249 6171
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 1394 6060 1400 6112
rect 1452 6060 1458 6112
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 4540 6100 4568 6208
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8895 6208 8953 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 10612 6236 10640 6267
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 14568 6313 14596 6344
rect 15562 6332 15568 6384
rect 15620 6332 15626 6384
rect 16669 6375 16727 6381
rect 16669 6341 16681 6375
rect 16715 6372 16727 6375
rect 16758 6372 16764 6384
rect 16715 6344 16764 6372
rect 16715 6341 16727 6344
rect 16669 6335 16727 6341
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 17034 6332 17040 6384
rect 17092 6332 17098 6384
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11664 6276 11897 6304
rect 11664 6264 11670 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16356 6276 16865 6304
rect 16356 6264 16362 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6304 17003 6307
rect 17052 6304 17080 6332
rect 17144 6313 17172 6412
rect 18782 6400 18788 6452
rect 18840 6440 18846 6452
rect 18877 6443 18935 6449
rect 18877 6440 18889 6443
rect 18840 6412 18889 6440
rect 18840 6400 18846 6412
rect 18877 6409 18889 6412
rect 18923 6409 18935 6443
rect 18877 6403 18935 6409
rect 17402 6332 17408 6384
rect 17460 6332 17466 6384
rect 18414 6332 18420 6384
rect 18472 6332 18478 6384
rect 16991 6276 17080 6304
rect 17129 6307 17187 6313
rect 16991 6273 17003 6276
rect 16945 6267 17003 6273
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 9364 6208 10640 6236
rect 9364 6196 9370 6208
rect 11698 6196 11704 6248
rect 11756 6196 11762 6248
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6236 12035 6239
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 12023 6208 12173 6236
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12802 6196 12808 6248
rect 12860 6196 12866 6248
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15856 6236 15884 6264
rect 18138 6236 18144 6248
rect 14875 6208 15884 6236
rect 15948 6208 18144 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 11808 6168 11836 6196
rect 15948 6168 15976 6208
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 11808 6140 12434 6168
rect 2188 6072 4568 6100
rect 2188 6060 2194 6072
rect 4614 6060 4620 6112
rect 4672 6060 4678 6112
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9585 6103 9643 6109
rect 9585 6100 9597 6103
rect 9272 6072 9597 6100
rect 9272 6060 9278 6072
rect 9585 6069 9597 6072
rect 9631 6069 9643 6103
rect 9585 6063 9643 6069
rect 9674 6060 9680 6112
rect 9732 6060 9738 6112
rect 10686 6060 10692 6112
rect 10744 6060 10750 6112
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 12406 6100 12434 6140
rect 15856 6140 15976 6168
rect 15856 6100 15884 6140
rect 16206 6128 16212 6180
rect 16264 6168 16270 6180
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 16264 6140 16313 6168
rect 16264 6128 16270 6140
rect 16301 6137 16313 6140
rect 16347 6168 16359 6171
rect 16850 6168 16856 6180
rect 16347 6140 16856 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 12406 6072 15884 6100
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 17862 6100 17868 6112
rect 15988 6072 17868 6100
rect 15988 6060 15994 6072
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 1104 6010 19228 6032
rect 1104 5958 3215 6010
rect 3267 5958 3279 6010
rect 3331 5958 3343 6010
rect 3395 5958 3407 6010
rect 3459 5958 3471 6010
rect 3523 5958 7746 6010
rect 7798 5958 7810 6010
rect 7862 5958 7874 6010
rect 7926 5958 7938 6010
rect 7990 5958 8002 6010
rect 8054 5958 12277 6010
rect 12329 5958 12341 6010
rect 12393 5958 12405 6010
rect 12457 5958 12469 6010
rect 12521 5958 12533 6010
rect 12585 5958 16808 6010
rect 16860 5958 16872 6010
rect 16924 5958 16936 6010
rect 16988 5958 17000 6010
rect 17052 5958 17064 6010
rect 17116 5958 19228 6010
rect 1104 5936 19228 5958
rect 1394 5856 1400 5908
rect 1452 5856 1458 5908
rect 2222 5856 2228 5908
rect 2280 5896 2286 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 2280 5868 2329 5896
rect 2280 5856 2286 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 2317 5859 2375 5865
rect 5368 5868 8217 5896
rect 1412 5692 1440 5856
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 2648 5732 2789 5760
rect 2648 5720 2654 5732
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 4246 5760 4252 5772
rect 2915 5732 4252 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 5368 5769 5396 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 9214 5896 9220 5908
rect 8205 5859 8263 5865
rect 8588 5868 9220 5896
rect 7377 5831 7435 5837
rect 7377 5797 7389 5831
rect 7423 5797 7435 5831
rect 7377 5791 7435 5797
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 5353 5763 5411 5769
rect 5353 5760 5365 5763
rect 4479 5732 5365 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 5353 5729 5365 5732
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 5905 5763 5963 5769
rect 5905 5760 5917 5763
rect 5583 5732 5917 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5905 5729 5917 5732
rect 5951 5729 5963 5763
rect 7392 5760 7420 5791
rect 8481 5763 8539 5769
rect 7392 5732 8432 5760
rect 5905 5723 5963 5729
rect 1489 5695 1547 5701
rect 1489 5692 1501 5695
rect 1412 5664 1501 5692
rect 1489 5661 1501 5664
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2685 5695 2743 5701
rect 2271 5664 2636 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 2498 5516 2504 5568
rect 2556 5516 2562 5568
rect 2608 5556 2636 5664
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2700 5624 2728 5655
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4614 5692 4620 5704
rect 4571 5664 4620 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 3786 5624 3792 5636
rect 2700 5596 3792 5624
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 5092 5624 5120 5655
rect 5166 5652 5172 5704
rect 5224 5652 5230 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5629 5695 5687 5701
rect 5629 5692 5641 5695
rect 5368 5664 5641 5692
rect 5368 5636 5396 5664
rect 5629 5661 5641 5664
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8404 5692 8432 5732
rect 8481 5729 8493 5763
rect 8527 5760 8539 5763
rect 8588 5760 8616 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9490 5856 9496 5908
rect 9548 5856 9554 5908
rect 9940 5899 9998 5905
rect 9940 5865 9952 5899
rect 9986 5896 9998 5899
rect 11514 5896 11520 5908
rect 9986 5868 11520 5896
rect 9986 5865 9998 5868
rect 9940 5859 9998 5865
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 12989 5899 13047 5905
rect 12989 5896 13001 5899
rect 12860 5868 13001 5896
rect 12860 5856 12866 5868
rect 12989 5865 13001 5868
rect 13035 5865 13047 5899
rect 12989 5859 13047 5865
rect 16666 5856 16672 5908
rect 16724 5856 16730 5908
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 17402 5896 17408 5908
rect 17083 5868 17408 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 18414 5896 18420 5908
rect 18371 5868 18420 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 11425 5831 11483 5837
rect 8812 5800 9444 5828
rect 8812 5788 8818 5800
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8527 5732 8616 5760
rect 8680 5732 9321 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8573 5695 8631 5701
rect 8404 5686 8524 5692
rect 8573 5686 8585 5695
rect 8404 5664 8585 5686
rect 8113 5655 8171 5661
rect 8496 5661 8585 5664
rect 8619 5694 8631 5695
rect 8680 5694 8708 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 8619 5666 8708 5694
rect 9125 5695 9183 5701
rect 8619 5661 8631 5666
rect 8496 5658 8631 5661
rect 8573 5655 8631 5658
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9214 5692 9220 5704
rect 9171 5664 9220 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 5092 5596 5212 5624
rect 2682 5556 2688 5568
rect 2608 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 4890 5516 4896 5568
rect 4948 5516 4954 5568
rect 5184 5556 5212 5596
rect 5350 5584 5356 5636
rect 5408 5584 5414 5636
rect 6914 5584 6920 5636
rect 6972 5584 6978 5636
rect 8128 5624 8156 5655
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9416 5701 9444 5800
rect 11425 5797 11437 5831
rect 11471 5828 11483 5831
rect 11882 5828 11888 5840
rect 11471 5800 11888 5828
rect 11471 5797 11483 5800
rect 11425 5791 11483 5797
rect 11882 5788 11888 5800
rect 11940 5828 11946 5840
rect 15841 5831 15899 5837
rect 11940 5800 13400 5828
rect 11940 5788 11946 5800
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10962 5760 10968 5772
rect 9723 5732 10968 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 13372 5769 13400 5800
rect 15841 5797 15853 5831
rect 15887 5828 15899 5831
rect 16022 5828 16028 5840
rect 15887 5800 16028 5828
rect 15887 5797 15899 5800
rect 15841 5791 15899 5797
rect 16022 5788 16028 5800
rect 16080 5828 16086 5840
rect 16684 5828 16712 5856
rect 16080 5800 16436 5828
rect 16684 5800 16804 5828
rect 16080 5788 16086 5800
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 11756 5732 12449 5760
rect 11756 5720 11762 5732
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 16298 5720 16304 5772
rect 16356 5720 16362 5772
rect 16408 5760 16436 5800
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 16408 5732 16681 5760
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12618 5692 12624 5704
rect 12575 5664 12624 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 8941 5627 8999 5633
rect 8941 5624 8953 5627
rect 8128 5596 8953 5624
rect 8941 5593 8953 5596
rect 8987 5593 8999 5627
rect 8941 5587 8999 5593
rect 10686 5584 10692 5636
rect 10744 5584 10750 5636
rect 13188 5624 13216 5655
rect 16206 5652 16212 5704
rect 16264 5701 16270 5704
rect 16776 5701 16804 5800
rect 16264 5692 16274 5701
rect 16761 5695 16819 5701
rect 16264 5664 16309 5692
rect 16264 5655 16274 5664
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 16264 5652 16270 5655
rect 17862 5652 17868 5704
rect 17920 5692 17926 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 17920 5664 18429 5692
rect 17920 5652 17926 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 12406 5596 13216 5624
rect 7469 5559 7527 5565
rect 7469 5556 7481 5559
rect 5184 5528 7481 5556
rect 7469 5525 7481 5528
rect 7515 5525 7527 5559
rect 7469 5519 7527 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12032 5528 12265 5556
rect 12032 5516 12038 5528
rect 12253 5525 12265 5528
rect 12299 5556 12311 5559
rect 12406 5556 12434 5596
rect 12299 5528 12434 5556
rect 12299 5525 12311 5528
rect 12253 5519 12311 5525
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12676 5528 12909 5556
rect 12676 5516 12682 5528
rect 12897 5525 12909 5528
rect 12943 5525 12955 5559
rect 12897 5519 12955 5525
rect 1104 5466 19228 5488
rect 1104 5414 3875 5466
rect 3927 5414 3939 5466
rect 3991 5414 4003 5466
rect 4055 5414 4067 5466
rect 4119 5414 4131 5466
rect 4183 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 8534 5466
rect 8586 5414 8598 5466
rect 8650 5414 8662 5466
rect 8714 5414 12937 5466
rect 12989 5414 13001 5466
rect 13053 5414 13065 5466
rect 13117 5414 13129 5466
rect 13181 5414 13193 5466
rect 13245 5414 17468 5466
rect 17520 5414 17532 5466
rect 17584 5414 17596 5466
rect 17648 5414 17660 5466
rect 17712 5414 17724 5466
rect 17776 5414 19228 5466
rect 1104 5392 19228 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 3016 5324 3157 5352
rect 3016 5312 3022 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 4890 5352 4896 5364
rect 3145 5315 3203 5321
rect 4724 5324 4896 5352
rect 4724 5293 4752 5324
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 6914 5352 6920 5364
rect 6779 5324 6920 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 9582 5352 9588 5364
rect 9232 5324 9588 5352
rect 4709 5287 4767 5293
rect 4709 5253 4721 5287
rect 4755 5253 4767 5287
rect 4709 5247 4767 5253
rect 5718 5244 5724 5296
rect 5776 5244 5782 5296
rect 9232 5293 9260 5324
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10689 5355 10747 5361
rect 10689 5321 10701 5355
rect 10735 5352 10747 5355
rect 11606 5352 11612 5364
rect 10735 5324 11612 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 14090 5352 14096 5364
rect 14047 5324 14096 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 14642 5312 14648 5364
rect 14700 5312 14706 5364
rect 15933 5355 15991 5361
rect 15933 5321 15945 5355
rect 15979 5352 15991 5355
rect 16298 5352 16304 5364
rect 15979 5324 16304 5352
rect 15979 5321 15991 5324
rect 15933 5315 15991 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 9217 5287 9275 5293
rect 7024 5256 8984 5284
rect 7024 5228 7052 5256
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 6641 5219 6699 5225
rect 3375 5188 4292 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 4264 5160 4292 5188
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 3605 5151 3663 5157
rect 3605 5148 3617 5151
rect 3559 5120 3617 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3605 5117 3617 5120
rect 3651 5117 3663 5151
rect 3605 5111 3663 5117
rect 4154 5108 4160 5160
rect 4212 5108 4218 5160
rect 4246 5108 4252 5160
rect 4304 5108 4310 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 5350 5148 5356 5160
rect 4479 5120 5356 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 1762 5040 1768 5092
rect 1820 5080 1826 5092
rect 2314 5080 2320 5092
rect 1820 5052 2320 5080
rect 1820 5040 1826 5052
rect 2314 5040 2320 5052
rect 2372 5080 2378 5092
rect 4448 5080 4476 5111
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 6656 5148 6684 5179
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 8956 5225 8984 5256
rect 9217 5253 9229 5287
rect 9263 5253 9275 5287
rect 9217 5247 9275 5253
rect 9674 5244 9680 5296
rect 9732 5244 9738 5296
rect 12529 5287 12587 5293
rect 10980 5256 12296 5284
rect 10980 5228 11008 5256
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 8941 5219 8999 5225
rect 8435 5188 8892 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 5500 5120 8585 5148
rect 5500 5108 5506 5120
rect 8573 5117 8585 5120
rect 8619 5148 8631 5151
rect 8754 5148 8760 5160
rect 8619 5120 8760 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8864 5148 8892 5188
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 10962 5176 10968 5228
rect 11020 5176 11026 5228
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 12268 5225 12296 5256
rect 12529 5253 12541 5287
rect 12575 5284 12587 5287
rect 12618 5284 12624 5296
rect 12575 5256 12624 5284
rect 12575 5253 12587 5256
rect 12529 5247 12587 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 13262 5244 13268 5296
rect 13320 5244 13326 5296
rect 14660 5284 14688 5312
rect 14200 5256 14688 5284
rect 14200 5225 14228 5256
rect 15102 5244 15108 5296
rect 15160 5244 15166 5296
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 9306 5148 9312 5160
rect 8864 5120 9312 5148
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5148 11575 5151
rect 11698 5148 11704 5160
rect 11563 5120 11704 5148
rect 11563 5117 11575 5120
rect 11517 5111 11575 5117
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 11974 5108 11980 5160
rect 12032 5108 12038 5160
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5148 14519 5151
rect 14918 5148 14924 5160
rect 14507 5120 14924 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 2372 5052 4476 5080
rect 2372 5040 2378 5052
rect 6178 4972 6184 5024
rect 6236 4972 6242 5024
rect 1104 4922 19228 4944
rect 1104 4870 3215 4922
rect 3267 4870 3279 4922
rect 3331 4870 3343 4922
rect 3395 4870 3407 4922
rect 3459 4870 3471 4922
rect 3523 4870 7746 4922
rect 7798 4870 7810 4922
rect 7862 4870 7874 4922
rect 7926 4870 7938 4922
rect 7990 4870 8002 4922
rect 8054 4870 12277 4922
rect 12329 4870 12341 4922
rect 12393 4870 12405 4922
rect 12457 4870 12469 4922
rect 12521 4870 12533 4922
rect 12585 4870 16808 4922
rect 16860 4870 16872 4922
rect 16924 4870 16936 4922
rect 16988 4870 17000 4922
rect 17052 4870 17064 4922
rect 17116 4870 19228 4922
rect 1104 4848 19228 4870
rect 3786 4768 3792 4820
rect 3844 4768 3850 4820
rect 4154 4768 4160 4820
rect 4212 4768 4218 4820
rect 5718 4768 5724 4820
rect 5776 4768 5782 4820
rect 6178 4768 6184 4820
rect 6236 4768 6242 4820
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9674 4808 9680 4820
rect 9539 4780 9680 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 13320 4780 13369 4808
rect 13320 4768 13326 4780
rect 13357 4777 13369 4780
rect 13403 4777 13415 4811
rect 13357 4771 13415 4777
rect 15102 4768 15108 4820
rect 15160 4768 15166 4820
rect 3513 4743 3571 4749
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 4172 4740 4200 4768
rect 3559 4712 4200 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 1762 4632 1768 4684
rect 1820 4632 1826 4684
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4672 2099 4675
rect 2498 4672 2504 4684
rect 2087 4644 2504 4672
rect 2087 4641 2099 4644
rect 2041 4635 2099 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 4172 4613 4200 4712
rect 4246 4632 4252 4684
rect 4304 4672 4310 4684
rect 6196 4672 6224 4768
rect 4304 4644 6224 4672
rect 4304 4632 4310 4644
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5500 4576 5825 4604
rect 5500 4564 5506 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8812 4576 9413 4604
rect 8812 4564 8818 4576
rect 9401 4573 9413 4576
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 12768 4576 13277 4604
rect 12768 4564 12774 4576
rect 13265 4573 13277 4576
rect 13311 4604 13323 4607
rect 14918 4604 14924 4616
rect 13311 4576 14924 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 14918 4564 14924 4576
rect 14976 4604 14982 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 14976 4576 15025 4604
rect 14976 4564 14982 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 2774 4496 2780 4548
rect 2832 4496 2838 4548
rect 1104 4378 19228 4400
rect 1104 4326 3875 4378
rect 3927 4326 3939 4378
rect 3991 4326 4003 4378
rect 4055 4326 4067 4378
rect 4119 4326 4131 4378
rect 4183 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 8534 4378
rect 8586 4326 8598 4378
rect 8650 4326 8662 4378
rect 8714 4326 12937 4378
rect 12989 4326 13001 4378
rect 13053 4326 13065 4378
rect 13117 4326 13129 4378
rect 13181 4326 13193 4378
rect 13245 4326 17468 4378
rect 17520 4326 17532 4378
rect 17584 4326 17596 4378
rect 17648 4326 17660 4378
rect 17712 4326 17724 4378
rect 17776 4326 19228 4378
rect 1104 4304 19228 4326
rect 2774 4224 2780 4276
rect 2832 4224 2838 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14976 4236 15025 4264
rect 14976 4224 14982 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 15286 4156 15292 4208
rect 15344 4156 15350 4208
rect 2682 4088 2688 4140
rect 2740 4088 2746 4140
rect 1104 3834 19228 3856
rect 1104 3782 3215 3834
rect 3267 3782 3279 3834
rect 3331 3782 3343 3834
rect 3395 3782 3407 3834
rect 3459 3782 3471 3834
rect 3523 3782 7746 3834
rect 7798 3782 7810 3834
rect 7862 3782 7874 3834
rect 7926 3782 7938 3834
rect 7990 3782 8002 3834
rect 8054 3782 12277 3834
rect 12329 3782 12341 3834
rect 12393 3782 12405 3834
rect 12457 3782 12469 3834
rect 12521 3782 12533 3834
rect 12585 3782 16808 3834
rect 16860 3782 16872 3834
rect 16924 3782 16936 3834
rect 16988 3782 17000 3834
rect 17052 3782 17064 3834
rect 17116 3782 19228 3834
rect 1104 3760 19228 3782
rect 1104 3290 19228 3312
rect 1104 3238 3875 3290
rect 3927 3238 3939 3290
rect 3991 3238 4003 3290
rect 4055 3238 4067 3290
rect 4119 3238 4131 3290
rect 4183 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 8534 3290
rect 8586 3238 8598 3290
rect 8650 3238 8662 3290
rect 8714 3238 12937 3290
rect 12989 3238 13001 3290
rect 13053 3238 13065 3290
rect 13117 3238 13129 3290
rect 13181 3238 13193 3290
rect 13245 3238 17468 3290
rect 17520 3238 17532 3290
rect 17584 3238 17596 3290
rect 17648 3238 17660 3290
rect 17712 3238 17724 3290
rect 17776 3238 19228 3290
rect 1104 3216 19228 3238
rect 1104 2746 19228 2768
rect 1104 2694 3215 2746
rect 3267 2694 3279 2746
rect 3331 2694 3343 2746
rect 3395 2694 3407 2746
rect 3459 2694 3471 2746
rect 3523 2694 7746 2746
rect 7798 2694 7810 2746
rect 7862 2694 7874 2746
rect 7926 2694 7938 2746
rect 7990 2694 8002 2746
rect 8054 2694 12277 2746
rect 12329 2694 12341 2746
rect 12393 2694 12405 2746
rect 12457 2694 12469 2746
rect 12521 2694 12533 2746
rect 12585 2694 16808 2746
rect 16860 2694 16872 2746
rect 16924 2694 16936 2746
rect 16988 2694 17000 2746
rect 17052 2694 17064 2746
rect 17116 2694 19228 2746
rect 1104 2672 19228 2694
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 15344 2604 15485 2632
rect 15344 2592 15350 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 1104 2202 19228 2224
rect 1104 2150 3875 2202
rect 3927 2150 3939 2202
rect 3991 2150 4003 2202
rect 4055 2150 4067 2202
rect 4119 2150 4131 2202
rect 4183 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 8534 2202
rect 8586 2150 8598 2202
rect 8650 2150 8662 2202
rect 8714 2150 12937 2202
rect 12989 2150 13001 2202
rect 13053 2150 13065 2202
rect 13117 2150 13129 2202
rect 13181 2150 13193 2202
rect 13245 2150 17468 2202
rect 17520 2150 17532 2202
rect 17584 2150 17596 2202
rect 17648 2150 17660 2202
rect 17712 2150 17724 2202
rect 17776 2150 19228 2202
rect 1104 2128 19228 2150
<< via1 >>
rect 16580 20340 16632 20392
rect 17500 20340 17552 20392
rect 3215 20102 3267 20154
rect 3279 20102 3331 20154
rect 3343 20102 3395 20154
rect 3407 20102 3459 20154
rect 3471 20102 3523 20154
rect 7746 20102 7798 20154
rect 7810 20102 7862 20154
rect 7874 20102 7926 20154
rect 7938 20102 7990 20154
rect 8002 20102 8054 20154
rect 12277 20102 12329 20154
rect 12341 20102 12393 20154
rect 12405 20102 12457 20154
rect 12469 20102 12521 20154
rect 12533 20102 12585 20154
rect 16808 20102 16860 20154
rect 16872 20102 16924 20154
rect 16936 20102 16988 20154
rect 17000 20102 17052 20154
rect 17064 20102 17116 20154
rect 3148 20000 3200 20052
rect 6552 20000 6604 20052
rect 13820 20000 13872 20052
rect 17868 20000 17920 20052
rect 2964 19932 3016 19984
rect 9220 19932 9272 19984
rect 1584 19796 1636 19848
rect 2136 19796 2188 19848
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 2780 19796 2832 19805
rect 3056 19796 3108 19848
rect 3792 19796 3844 19848
rect 4344 19796 4396 19848
rect 4896 19796 4948 19848
rect 5540 19796 5592 19848
rect 6000 19796 6052 19848
rect 13176 19864 13228 19916
rect 7104 19796 7156 19848
rect 7656 19796 7708 19848
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 8760 19796 8812 19848
rect 9312 19796 9364 19848
rect 9864 19796 9916 19848
rect 10416 19796 10468 19848
rect 11060 19839 11112 19848
rect 11060 19805 11069 19839
rect 11069 19805 11103 19839
rect 11103 19805 11112 19839
rect 11060 19796 11112 19805
rect 11520 19796 11572 19848
rect 12072 19796 12124 19848
rect 12624 19796 12676 19848
rect 14280 19796 14332 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 15752 19932 15804 19984
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15384 19796 15436 19848
rect 15936 19796 15988 19848
rect 16580 19796 16632 19848
rect 17960 19932 18012 19984
rect 17224 19864 17276 19916
rect 17592 19864 17644 19916
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 2136 19660 2188 19712
rect 3516 19703 3568 19712
rect 3516 19669 3525 19703
rect 3525 19669 3559 19703
rect 3559 19669 3568 19703
rect 3516 19660 3568 19669
rect 4528 19660 4580 19712
rect 4620 19703 4672 19712
rect 4620 19669 4629 19703
rect 4629 19669 4663 19703
rect 4663 19669 4672 19703
rect 4620 19660 4672 19669
rect 4988 19703 5040 19712
rect 4988 19669 4997 19703
rect 4997 19669 5031 19703
rect 5031 19669 5040 19703
rect 4988 19660 5040 19669
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 6552 19660 6604 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 7380 19660 7432 19712
rect 8944 19703 8996 19712
rect 8944 19669 8953 19703
rect 8953 19669 8987 19703
rect 8987 19669 8996 19703
rect 8944 19660 8996 19669
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 10140 19703 10192 19712
rect 10140 19669 10149 19703
rect 10149 19669 10183 19703
rect 10183 19669 10192 19703
rect 10140 19660 10192 19669
rect 10784 19660 10836 19712
rect 11244 19703 11296 19712
rect 11244 19669 11253 19703
rect 11253 19669 11287 19703
rect 11287 19669 11296 19703
rect 11244 19660 11296 19669
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 11888 19660 11940 19712
rect 13452 19660 13504 19712
rect 13636 19660 13688 19712
rect 13728 19703 13780 19712
rect 13728 19669 13737 19703
rect 13737 19669 13771 19703
rect 13771 19669 13780 19703
rect 13728 19660 13780 19669
rect 14004 19660 14056 19712
rect 14188 19703 14240 19712
rect 14188 19669 14197 19703
rect 14197 19669 14231 19703
rect 14231 19669 14240 19703
rect 14188 19660 14240 19669
rect 15108 19703 15160 19712
rect 15108 19669 15117 19703
rect 15117 19669 15151 19703
rect 15151 19669 15160 19703
rect 15108 19660 15160 19669
rect 15384 19660 15436 19712
rect 15476 19660 15528 19712
rect 16212 19703 16264 19712
rect 16212 19669 16221 19703
rect 16221 19669 16255 19703
rect 16255 19669 16264 19703
rect 16212 19660 16264 19669
rect 16672 19703 16724 19712
rect 16672 19669 16681 19703
rect 16681 19669 16715 19703
rect 16715 19669 16724 19703
rect 16672 19660 16724 19669
rect 17500 19839 17552 19848
rect 17500 19805 17509 19839
rect 17509 19805 17543 19839
rect 17543 19805 17552 19839
rect 17500 19796 17552 19805
rect 18144 19796 18196 19848
rect 18696 19796 18748 19848
rect 17316 19660 17368 19712
rect 17408 19660 17460 19712
rect 17684 19660 17736 19712
rect 18236 19703 18288 19712
rect 18236 19669 18245 19703
rect 18245 19669 18279 19703
rect 18279 19669 18288 19703
rect 18236 19660 18288 19669
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 3875 19558 3927 19610
rect 3939 19558 3991 19610
rect 4003 19558 4055 19610
rect 4067 19558 4119 19610
rect 4131 19558 4183 19610
rect 8406 19558 8458 19610
rect 8470 19558 8522 19610
rect 8534 19558 8586 19610
rect 8598 19558 8650 19610
rect 8662 19558 8714 19610
rect 12937 19558 12989 19610
rect 13001 19558 13053 19610
rect 13065 19558 13117 19610
rect 13129 19558 13181 19610
rect 13193 19558 13245 19610
rect 17468 19558 17520 19610
rect 17532 19558 17584 19610
rect 17596 19558 17648 19610
rect 17660 19558 17712 19610
rect 17724 19558 17776 19610
rect 9036 19388 9088 19440
rect 2780 19320 2832 19372
rect 3884 19320 3936 19372
rect 2872 19252 2924 19304
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 2596 19184 2648 19236
rect 3976 19252 4028 19304
rect 4252 19320 4304 19372
rect 5816 19320 5868 19372
rect 6828 19320 6880 19372
rect 10140 19456 10192 19508
rect 10324 19456 10376 19508
rect 9772 19320 9824 19372
rect 10140 19320 10192 19372
rect 14372 19456 14424 19508
rect 14556 19456 14608 19508
rect 16672 19456 16724 19508
rect 11060 19388 11112 19440
rect 11336 19320 11388 19372
rect 13636 19388 13688 19440
rect 17408 19388 17460 19440
rect 4344 19252 4396 19304
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 9680 19252 9732 19304
rect 11152 19252 11204 19304
rect 12624 19295 12676 19304
rect 12624 19261 12633 19295
rect 12633 19261 12667 19295
rect 12667 19261 12676 19295
rect 12624 19252 12676 19261
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 2780 19159 2832 19168
rect 2780 19125 2789 19159
rect 2789 19125 2823 19159
rect 2823 19125 2832 19159
rect 2780 19116 2832 19125
rect 3792 19116 3844 19168
rect 4436 19184 4488 19236
rect 4896 19116 4948 19168
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 10232 19159 10284 19168
rect 10232 19125 10241 19159
rect 10241 19125 10275 19159
rect 10275 19125 10284 19159
rect 10232 19116 10284 19125
rect 11612 19159 11664 19168
rect 11612 19125 11621 19159
rect 11621 19125 11655 19159
rect 11655 19125 11664 19159
rect 11612 19116 11664 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 15384 19116 15436 19168
rect 16304 19116 16356 19168
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 3215 19014 3267 19066
rect 3279 19014 3331 19066
rect 3343 19014 3395 19066
rect 3407 19014 3459 19066
rect 3471 19014 3523 19066
rect 7746 19014 7798 19066
rect 7810 19014 7862 19066
rect 7874 19014 7926 19066
rect 7938 19014 7990 19066
rect 8002 19014 8054 19066
rect 12277 19014 12329 19066
rect 12341 19014 12393 19066
rect 12405 19014 12457 19066
rect 12469 19014 12521 19066
rect 12533 19014 12585 19066
rect 16808 19014 16860 19066
rect 16872 19014 16924 19066
rect 16936 19014 16988 19066
rect 17000 19014 17052 19066
rect 17064 19014 17116 19066
rect 2688 18912 2740 18964
rect 3976 18912 4028 18964
rect 4712 18912 4764 18964
rect 7288 18912 7340 18964
rect 8852 18912 8904 18964
rect 9312 18912 9364 18964
rect 10140 18912 10192 18964
rect 10232 18912 10284 18964
rect 12624 18912 12676 18964
rect 3700 18844 3752 18896
rect 4436 18844 4488 18896
rect 5356 18819 5408 18828
rect 5356 18785 5365 18819
rect 5365 18785 5399 18819
rect 5399 18785 5408 18819
rect 5356 18776 5408 18785
rect 5540 18844 5592 18896
rect 6368 18844 6420 18896
rect 6184 18776 6236 18828
rect 6644 18819 6696 18828
rect 6644 18785 6653 18819
rect 6653 18785 6687 18819
rect 6687 18785 6696 18819
rect 6644 18776 6696 18785
rect 9772 18776 9824 18828
rect 10140 18776 10192 18828
rect 10968 18776 11020 18828
rect 13268 18819 13320 18828
rect 13268 18785 13277 18819
rect 13277 18785 13311 18819
rect 13311 18785 13320 18819
rect 13268 18776 13320 18785
rect 13728 18776 13780 18828
rect 14188 18776 14240 18828
rect 16304 18912 16356 18964
rect 17408 18955 17460 18964
rect 17408 18921 17417 18955
rect 17417 18921 17451 18955
rect 17451 18921 17460 18955
rect 17408 18912 17460 18921
rect 16580 18844 16632 18896
rect 3148 18708 3200 18760
rect 4436 18708 4488 18760
rect 4896 18708 4948 18760
rect 1768 18572 1820 18624
rect 2596 18640 2648 18692
rect 3884 18640 3936 18692
rect 6000 18640 6052 18692
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 11612 18708 11664 18760
rect 9404 18640 9456 18692
rect 14556 18708 14608 18760
rect 13636 18640 13688 18692
rect 16764 18776 16816 18828
rect 18512 18844 18564 18896
rect 16672 18708 16724 18760
rect 18420 18776 18472 18828
rect 15200 18683 15252 18692
rect 15200 18649 15209 18683
rect 15209 18649 15243 18683
rect 15243 18649 15252 18683
rect 15200 18640 15252 18649
rect 2780 18572 2832 18624
rect 8484 18572 8536 18624
rect 10416 18572 10468 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 13544 18572 13596 18624
rect 16580 18572 16632 18624
rect 3875 18470 3927 18522
rect 3939 18470 3991 18522
rect 4003 18470 4055 18522
rect 4067 18470 4119 18522
rect 4131 18470 4183 18522
rect 8406 18470 8458 18522
rect 8470 18470 8522 18522
rect 8534 18470 8586 18522
rect 8598 18470 8650 18522
rect 8662 18470 8714 18522
rect 12937 18470 12989 18522
rect 13001 18470 13053 18522
rect 13065 18470 13117 18522
rect 13129 18470 13181 18522
rect 13193 18470 13245 18522
rect 17468 18470 17520 18522
rect 17532 18470 17584 18522
rect 17596 18470 17648 18522
rect 17660 18470 17712 18522
rect 17724 18470 17776 18522
rect 3792 18368 3844 18420
rect 4344 18368 4396 18420
rect 5540 18368 5592 18420
rect 5816 18368 5868 18420
rect 6644 18368 6696 18420
rect 9404 18368 9456 18420
rect 9680 18368 9732 18420
rect 9864 18368 9916 18420
rect 13728 18368 13780 18420
rect 15200 18368 15252 18420
rect 15292 18368 15344 18420
rect 1768 18232 1820 18284
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 4252 18300 4304 18352
rect 3148 18232 3200 18241
rect 3700 18232 3752 18284
rect 3792 18232 3844 18284
rect 2872 18164 2924 18216
rect 4436 18164 4488 18216
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 6920 18232 6972 18284
rect 5356 18164 5408 18216
rect 7564 18164 7616 18216
rect 4804 18028 4856 18080
rect 5908 18028 5960 18080
rect 8852 18232 8904 18284
rect 9312 18300 9364 18352
rect 9956 18232 10008 18284
rect 9036 18164 9088 18216
rect 9680 18096 9732 18148
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 12072 18300 12124 18352
rect 18512 18300 18564 18352
rect 10416 18207 10468 18216
rect 10416 18173 10425 18207
rect 10425 18173 10459 18207
rect 10459 18173 10468 18207
rect 10416 18164 10468 18173
rect 11060 18164 11112 18216
rect 11980 18164 12032 18216
rect 11152 18096 11204 18148
rect 16764 18164 16816 18216
rect 17960 18164 18012 18216
rect 15384 18096 15436 18148
rect 11336 18028 11388 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 15844 18028 15896 18080
rect 3215 17926 3267 17978
rect 3279 17926 3331 17978
rect 3343 17926 3395 17978
rect 3407 17926 3459 17978
rect 3471 17926 3523 17978
rect 7746 17926 7798 17978
rect 7810 17926 7862 17978
rect 7874 17926 7926 17978
rect 7938 17926 7990 17978
rect 8002 17926 8054 17978
rect 12277 17926 12329 17978
rect 12341 17926 12393 17978
rect 12405 17926 12457 17978
rect 12469 17926 12521 17978
rect 12533 17926 12585 17978
rect 16808 17926 16860 17978
rect 16872 17926 16924 17978
rect 16936 17926 16988 17978
rect 17000 17926 17052 17978
rect 17064 17926 17116 17978
rect 7564 17824 7616 17876
rect 10048 17824 10100 17876
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 12348 17688 12400 17740
rect 13268 17731 13320 17740
rect 13268 17697 13277 17731
rect 13277 17697 13311 17731
rect 13311 17697 13320 17731
rect 13268 17688 13320 17697
rect 16672 17688 16724 17740
rect 2872 17620 2924 17672
rect 3056 17620 3108 17672
rect 3792 17620 3844 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 15108 17620 15160 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 5724 17595 5776 17604
rect 5724 17561 5733 17595
rect 5733 17561 5767 17595
rect 5767 17561 5776 17595
rect 5724 17552 5776 17561
rect 6460 17552 6512 17604
rect 11152 17552 11204 17604
rect 17040 17595 17092 17604
rect 17040 17561 17049 17595
rect 17049 17561 17083 17595
rect 17083 17561 17092 17595
rect 17040 17552 17092 17561
rect 18052 17552 18104 17604
rect 12808 17484 12860 17536
rect 13728 17527 13780 17536
rect 13728 17493 13737 17527
rect 13737 17493 13771 17527
rect 13771 17493 13780 17527
rect 13728 17484 13780 17493
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 16120 17484 16172 17536
rect 3875 17382 3927 17434
rect 3939 17382 3991 17434
rect 4003 17382 4055 17434
rect 4067 17382 4119 17434
rect 4131 17382 4183 17434
rect 8406 17382 8458 17434
rect 8470 17382 8522 17434
rect 8534 17382 8586 17434
rect 8598 17382 8650 17434
rect 8662 17382 8714 17434
rect 12937 17382 12989 17434
rect 13001 17382 13053 17434
rect 13065 17382 13117 17434
rect 13129 17382 13181 17434
rect 13193 17382 13245 17434
rect 17468 17382 17520 17434
rect 17532 17382 17584 17434
rect 17596 17382 17648 17434
rect 17660 17382 17712 17434
rect 17724 17382 17776 17434
rect 2688 17280 2740 17332
rect 3148 17280 3200 17332
rect 940 17144 992 17196
rect 2044 17144 2096 17196
rect 4804 17280 4856 17332
rect 5080 17212 5132 17264
rect 2688 17076 2740 17128
rect 3056 17076 3108 17128
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 2872 16940 2924 16992
rect 4620 16983 4672 16992
rect 4620 16949 4629 16983
rect 4629 16949 4663 16983
rect 4663 16949 4672 16983
rect 4620 16940 4672 16949
rect 4896 16940 4948 16992
rect 5264 17076 5316 17128
rect 6552 17280 6604 17332
rect 11152 17280 11204 17332
rect 12348 17280 12400 17332
rect 12808 17280 12860 17332
rect 13728 17280 13780 17332
rect 5908 17193 5960 17196
rect 5908 17159 5917 17193
rect 5917 17159 5951 17193
rect 5951 17159 5960 17193
rect 5908 17144 5960 17159
rect 11336 17212 11388 17264
rect 5724 17008 5776 17060
rect 8300 17144 8352 17196
rect 15844 17280 15896 17332
rect 17040 17280 17092 17332
rect 18052 17280 18104 17332
rect 12808 17187 12860 17196
rect 8484 17119 8536 17128
rect 8484 17085 8493 17119
rect 8493 17085 8527 17119
rect 8527 17085 8536 17119
rect 8484 17076 8536 17085
rect 11980 17119 12032 17128
rect 11980 17085 11989 17119
rect 11989 17085 12023 17119
rect 12023 17085 12032 17119
rect 11980 17076 12032 17085
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 14004 17076 14056 17128
rect 16580 17144 16632 17196
rect 11060 17008 11112 17060
rect 14924 17008 14976 17060
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 5080 16940 5132 16992
rect 5908 16940 5960 16992
rect 6920 16940 6972 16992
rect 8116 16940 8168 16992
rect 13544 16940 13596 16992
rect 16580 17008 16632 17060
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 15844 16940 15896 16992
rect 17316 16940 17368 16992
rect 18144 16940 18196 16992
rect 3215 16838 3267 16890
rect 3279 16838 3331 16890
rect 3343 16838 3395 16890
rect 3407 16838 3459 16890
rect 3471 16838 3523 16890
rect 7746 16838 7798 16890
rect 7810 16838 7862 16890
rect 7874 16838 7926 16890
rect 7938 16838 7990 16890
rect 8002 16838 8054 16890
rect 12277 16838 12329 16890
rect 12341 16838 12393 16890
rect 12405 16838 12457 16890
rect 12469 16838 12521 16890
rect 12533 16838 12585 16890
rect 16808 16838 16860 16890
rect 16872 16838 16924 16890
rect 16936 16838 16988 16890
rect 17000 16838 17052 16890
rect 17064 16838 17116 16890
rect 6460 16736 6512 16788
rect 8484 16736 8536 16788
rect 8760 16736 8812 16788
rect 10140 16736 10192 16788
rect 10692 16779 10744 16788
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 4620 16600 4672 16652
rect 8116 16668 8168 16720
rect 8944 16600 8996 16652
rect 15108 16600 15160 16652
rect 16764 16736 16816 16788
rect 16028 16668 16080 16720
rect 3792 16575 3844 16584
rect 2228 16464 2280 16516
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 4528 16464 4580 16516
rect 8300 16532 8352 16584
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 16672 16600 16724 16652
rect 18512 16600 18564 16652
rect 12164 16507 12216 16516
rect 12164 16473 12173 16507
rect 12173 16473 12207 16507
rect 12207 16473 12216 16507
rect 12164 16464 12216 16473
rect 2780 16396 2832 16448
rect 3056 16396 3108 16448
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 6460 16396 6512 16448
rect 7380 16439 7432 16448
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 7380 16396 7432 16405
rect 7656 16396 7708 16448
rect 17316 16464 17368 16516
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 3875 16294 3927 16346
rect 3939 16294 3991 16346
rect 4003 16294 4055 16346
rect 4067 16294 4119 16346
rect 4131 16294 4183 16346
rect 8406 16294 8458 16346
rect 8470 16294 8522 16346
rect 8534 16294 8586 16346
rect 8598 16294 8650 16346
rect 8662 16294 8714 16346
rect 12937 16294 12989 16346
rect 13001 16294 13053 16346
rect 13065 16294 13117 16346
rect 13129 16294 13181 16346
rect 13193 16294 13245 16346
rect 17468 16294 17520 16346
rect 17532 16294 17584 16346
rect 17596 16294 17648 16346
rect 17660 16294 17712 16346
rect 17724 16294 17776 16346
rect 4528 16235 4580 16244
rect 4528 16201 4537 16235
rect 4537 16201 4571 16235
rect 4571 16201 4580 16235
rect 4528 16192 4580 16201
rect 1584 16124 1636 16176
rect 5540 16192 5592 16244
rect 6276 16192 6328 16244
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 8760 16192 8812 16244
rect 9496 16192 9548 16244
rect 9680 16192 9732 16244
rect 5264 16124 5316 16176
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 6368 16056 6420 16108
rect 6828 16124 6880 16176
rect 7472 16124 7524 16176
rect 7380 15988 7432 16040
rect 9864 16124 9916 16176
rect 12808 16192 12860 16244
rect 16580 16192 16632 16244
rect 16764 16192 16816 16244
rect 17316 16192 17368 16244
rect 18236 16192 18288 16244
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 12072 16124 12124 16176
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 6460 15920 6512 15972
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 14924 15988 14976 16040
rect 18512 16099 18564 16108
rect 18512 16065 18521 16099
rect 18521 16065 18555 16099
rect 18555 16065 18564 16099
rect 18512 16056 18564 16065
rect 18880 15988 18932 16040
rect 18144 15963 18196 15972
rect 18144 15929 18153 15963
rect 18153 15929 18187 15963
rect 18187 15929 18196 15963
rect 18144 15920 18196 15929
rect 4252 15852 4304 15904
rect 5080 15852 5132 15904
rect 11152 15852 11204 15904
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 16120 15852 16172 15904
rect 3215 15750 3267 15802
rect 3279 15750 3331 15802
rect 3343 15750 3395 15802
rect 3407 15750 3459 15802
rect 3471 15750 3523 15802
rect 7746 15750 7798 15802
rect 7810 15750 7862 15802
rect 7874 15750 7926 15802
rect 7938 15750 7990 15802
rect 8002 15750 8054 15802
rect 12277 15750 12329 15802
rect 12341 15750 12393 15802
rect 12405 15750 12457 15802
rect 12469 15750 12521 15802
rect 12533 15750 12585 15802
rect 16808 15750 16860 15802
rect 16872 15750 16924 15802
rect 16936 15750 16988 15802
rect 17000 15750 17052 15802
rect 17064 15750 17116 15802
rect 7472 15648 7524 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 12072 15648 12124 15700
rect 13820 15648 13872 15700
rect 2228 15555 2280 15564
rect 2228 15521 2237 15555
rect 2237 15521 2271 15555
rect 2271 15521 2280 15555
rect 2228 15512 2280 15521
rect 2780 15512 2832 15564
rect 3424 15512 3476 15564
rect 8116 15580 8168 15632
rect 8760 15580 8812 15632
rect 9956 15580 10008 15632
rect 10968 15580 11020 15632
rect 3148 15444 3200 15496
rect 6460 15444 6512 15496
rect 6920 15376 6972 15428
rect 8944 15444 8996 15496
rect 10784 15512 10836 15564
rect 13636 15512 13688 15564
rect 14464 15512 14516 15564
rect 15384 15444 15436 15496
rect 12440 15419 12492 15428
rect 12440 15385 12449 15419
rect 12449 15385 12483 15419
rect 12483 15385 12492 15419
rect 12440 15376 12492 15385
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 6276 15308 6328 15360
rect 11520 15308 11572 15360
rect 13912 15308 13964 15360
rect 14280 15308 14332 15360
rect 3875 15206 3927 15258
rect 3939 15206 3991 15258
rect 4003 15206 4055 15258
rect 4067 15206 4119 15258
rect 4131 15206 4183 15258
rect 8406 15206 8458 15258
rect 8470 15206 8522 15258
rect 8534 15206 8586 15258
rect 8598 15206 8650 15258
rect 8662 15206 8714 15258
rect 12937 15206 12989 15258
rect 13001 15206 13053 15258
rect 13065 15206 13117 15258
rect 13129 15206 13181 15258
rect 13193 15206 13245 15258
rect 17468 15206 17520 15258
rect 17532 15206 17584 15258
rect 17596 15206 17648 15258
rect 17660 15206 17712 15258
rect 17724 15206 17776 15258
rect 3148 15147 3200 15156
rect 3148 15113 3157 15147
rect 3157 15113 3191 15147
rect 3191 15113 3200 15147
rect 3148 15104 3200 15113
rect 7196 15104 7248 15156
rect 12440 15104 12492 15156
rect 13452 15104 13504 15156
rect 15752 15104 15804 15156
rect 2136 15036 2188 15088
rect 3424 15011 3476 15020
rect 3424 14977 3433 15011
rect 3433 14977 3467 15011
rect 3467 14977 3476 15011
rect 3424 14968 3476 14977
rect 3792 14968 3844 15020
rect 6920 14968 6972 15020
rect 10416 15036 10468 15088
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 13912 15011 13964 15020
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 14280 14968 14332 15020
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 2780 14832 2832 14884
rect 9864 14900 9916 14952
rect 11704 14900 11756 14952
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 15384 14900 15436 14952
rect 16028 14968 16080 15020
rect 17500 15011 17552 15020
rect 17500 14977 17509 15011
rect 17509 14977 17543 15011
rect 17543 14977 17552 15011
rect 17500 14968 17552 14977
rect 18236 14900 18288 14952
rect 16120 14832 16172 14884
rect 6460 14807 6512 14816
rect 6460 14773 6469 14807
rect 6469 14773 6503 14807
rect 6503 14773 6512 14807
rect 6460 14764 6512 14773
rect 7012 14764 7064 14816
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 10876 14764 10928 14816
rect 13544 14764 13596 14816
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 15936 14807 15988 14816
rect 15936 14773 15945 14807
rect 15945 14773 15979 14807
rect 15979 14773 15988 14807
rect 15936 14764 15988 14773
rect 16580 14764 16632 14816
rect 17868 14764 17920 14816
rect 3215 14662 3267 14714
rect 3279 14662 3331 14714
rect 3343 14662 3395 14714
rect 3407 14662 3459 14714
rect 3471 14662 3523 14714
rect 7746 14662 7798 14714
rect 7810 14662 7862 14714
rect 7874 14662 7926 14714
rect 7938 14662 7990 14714
rect 8002 14662 8054 14714
rect 12277 14662 12329 14714
rect 12341 14662 12393 14714
rect 12405 14662 12457 14714
rect 12469 14662 12521 14714
rect 12533 14662 12585 14714
rect 16808 14662 16860 14714
rect 16872 14662 16924 14714
rect 16936 14662 16988 14714
rect 17000 14662 17052 14714
rect 17064 14662 17116 14714
rect 1676 14560 1728 14612
rect 5540 14603 5592 14612
rect 5540 14569 5549 14603
rect 5549 14569 5583 14603
rect 5583 14569 5592 14603
rect 5540 14560 5592 14569
rect 6460 14560 6512 14612
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 9864 14560 9916 14612
rect 10508 14560 10560 14612
rect 10876 14560 10928 14612
rect 2136 14535 2188 14544
rect 2136 14501 2145 14535
rect 2145 14501 2179 14535
rect 2179 14501 2188 14535
rect 2136 14492 2188 14501
rect 2228 14424 2280 14476
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 3056 14424 3108 14476
rect 6736 14492 6788 14544
rect 7656 14492 7708 14544
rect 7104 14424 7156 14476
rect 10692 14424 10744 14476
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 3700 14288 3752 14340
rect 6276 14288 6328 14340
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 7472 14356 7524 14408
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 13544 14560 13596 14612
rect 13820 14560 13872 14612
rect 16948 14560 17000 14612
rect 17500 14560 17552 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 13636 14424 13688 14476
rect 14372 14424 14424 14476
rect 16672 14424 16724 14476
rect 7196 14288 7248 14340
rect 18512 14356 18564 14408
rect 10876 14288 10928 14340
rect 15292 14331 15344 14340
rect 15292 14297 15301 14331
rect 15301 14297 15335 14331
rect 15335 14297 15344 14331
rect 15292 14288 15344 14297
rect 15936 14288 15988 14340
rect 17316 14288 17368 14340
rect 4988 14220 5040 14272
rect 6552 14220 6604 14272
rect 9036 14220 9088 14272
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 11796 14263 11848 14272
rect 11796 14229 11805 14263
rect 11805 14229 11839 14263
rect 11839 14229 11848 14263
rect 11796 14220 11848 14229
rect 13268 14220 13320 14272
rect 16028 14220 16080 14272
rect 16304 14220 16356 14272
rect 18052 14220 18104 14272
rect 3875 14118 3927 14170
rect 3939 14118 3991 14170
rect 4003 14118 4055 14170
rect 4067 14118 4119 14170
rect 4131 14118 4183 14170
rect 8406 14118 8458 14170
rect 8470 14118 8522 14170
rect 8534 14118 8586 14170
rect 8598 14118 8650 14170
rect 8662 14118 8714 14170
rect 12937 14118 12989 14170
rect 13001 14118 13053 14170
rect 13065 14118 13117 14170
rect 13129 14118 13181 14170
rect 13193 14118 13245 14170
rect 17468 14118 17520 14170
rect 17532 14118 17584 14170
rect 17596 14118 17648 14170
rect 17660 14118 17712 14170
rect 17724 14118 17776 14170
rect 3056 14016 3108 14068
rect 4252 13948 4304 14000
rect 4896 13948 4948 14000
rect 6552 13948 6604 14000
rect 10876 14016 10928 14068
rect 11704 14016 11756 14068
rect 11796 14016 11848 14068
rect 13544 14016 13596 14068
rect 15292 14016 15344 14068
rect 18052 14016 18104 14068
rect 18512 14059 18564 14068
rect 18512 14025 18521 14059
rect 18521 14025 18555 14059
rect 18555 14025 18564 14059
rect 18512 14016 18564 14025
rect 9128 13948 9180 14000
rect 2228 13812 2280 13864
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 10968 13880 11020 13932
rect 6276 13812 6328 13864
rect 6368 13855 6420 13864
rect 6368 13821 6377 13855
rect 6377 13821 6411 13855
rect 6411 13821 6420 13855
rect 6368 13812 6420 13821
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15752 13880 15804 13932
rect 17868 13948 17920 14000
rect 18236 13880 18288 13932
rect 12808 13812 12860 13864
rect 13268 13812 13320 13864
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 3700 13744 3752 13796
rect 4252 13676 4304 13728
rect 15660 13744 15712 13796
rect 15844 13744 15896 13796
rect 16948 13812 17000 13864
rect 7012 13676 7064 13728
rect 8116 13719 8168 13728
rect 8116 13685 8125 13719
rect 8125 13685 8159 13719
rect 8159 13685 8168 13719
rect 8116 13676 8168 13685
rect 8760 13676 8812 13728
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 17040 13676 17092 13728
rect 17224 13676 17276 13728
rect 3215 13574 3267 13626
rect 3279 13574 3331 13626
rect 3343 13574 3395 13626
rect 3407 13574 3459 13626
rect 3471 13574 3523 13626
rect 7746 13574 7798 13626
rect 7810 13574 7862 13626
rect 7874 13574 7926 13626
rect 7938 13574 7990 13626
rect 8002 13574 8054 13626
rect 12277 13574 12329 13626
rect 12341 13574 12393 13626
rect 12405 13574 12457 13626
rect 12469 13574 12521 13626
rect 12533 13574 12585 13626
rect 16808 13574 16860 13626
rect 16872 13574 16924 13626
rect 16936 13574 16988 13626
rect 17000 13574 17052 13626
rect 17064 13574 17116 13626
rect 6368 13472 6420 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 12808 13472 12860 13524
rect 17316 13472 17368 13524
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 6184 13336 6236 13388
rect 7656 13404 7708 13456
rect 2044 13268 2096 13320
rect 5632 13268 5684 13320
rect 8116 13336 8168 13388
rect 10692 13336 10744 13388
rect 17868 13336 17920 13388
rect 9036 13268 9088 13320
rect 5264 13243 5316 13252
rect 5264 13209 5273 13243
rect 5273 13209 5307 13243
rect 5307 13209 5316 13243
rect 5264 13200 5316 13209
rect 10048 13268 10100 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 16580 13268 16632 13320
rect 11060 13243 11112 13252
rect 11060 13209 11069 13243
rect 11069 13209 11103 13243
rect 11103 13209 11112 13243
rect 11060 13200 11112 13209
rect 11796 13200 11848 13252
rect 4896 13132 4948 13184
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 8944 13132 8996 13184
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 3875 13030 3927 13082
rect 3939 13030 3991 13082
rect 4003 13030 4055 13082
rect 4067 13030 4119 13082
rect 4131 13030 4183 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 8534 13030 8586 13082
rect 8598 13030 8650 13082
rect 8662 13030 8714 13082
rect 12937 13030 12989 13082
rect 13001 13030 13053 13082
rect 13065 13030 13117 13082
rect 13129 13030 13181 13082
rect 13193 13030 13245 13082
rect 17468 13030 17520 13082
rect 17532 13030 17584 13082
rect 17596 13030 17648 13082
rect 17660 13030 17712 13082
rect 17724 13030 17776 13082
rect 4896 12928 4948 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 7472 12971 7524 12980
rect 7472 12937 7481 12971
rect 7481 12937 7515 12971
rect 7515 12937 7524 12971
rect 7472 12928 7524 12937
rect 4252 12860 4304 12912
rect 2688 12792 2740 12844
rect 7656 12835 7708 12844
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 8116 12928 8168 12980
rect 10232 12928 10284 12980
rect 11060 12971 11112 12980
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 11152 12928 11204 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 14372 12928 14424 12980
rect 15476 12928 15528 12980
rect 18236 12928 18288 12980
rect 8300 12860 8352 12912
rect 8944 12860 8996 12912
rect 11244 12792 11296 12844
rect 12624 12860 12676 12912
rect 18420 12860 18472 12912
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16672 12792 16724 12844
rect 6368 12656 6420 12708
rect 8944 12724 8996 12776
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 16672 12656 16724 12708
rect 3884 12631 3936 12640
rect 3884 12597 3893 12631
rect 3893 12597 3927 12631
rect 3927 12597 3936 12631
rect 3884 12588 3936 12597
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 18052 12588 18104 12640
rect 3215 12486 3267 12538
rect 3279 12486 3331 12538
rect 3343 12486 3395 12538
rect 3407 12486 3459 12538
rect 3471 12486 3523 12538
rect 7746 12486 7798 12538
rect 7810 12486 7862 12538
rect 7874 12486 7926 12538
rect 7938 12486 7990 12538
rect 8002 12486 8054 12538
rect 12277 12486 12329 12538
rect 12341 12486 12393 12538
rect 12405 12486 12457 12538
rect 12469 12486 12521 12538
rect 12533 12486 12585 12538
rect 16808 12486 16860 12538
rect 16872 12486 16924 12538
rect 16936 12486 16988 12538
rect 17000 12486 17052 12538
rect 17064 12486 17116 12538
rect 5632 12427 5684 12436
rect 5632 12393 5641 12427
rect 5641 12393 5675 12427
rect 5675 12393 5684 12427
rect 5632 12384 5684 12393
rect 7656 12384 7708 12436
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 3884 12291 3936 12300
rect 1400 12248 1452 12257
rect 3884 12257 3893 12291
rect 3893 12257 3927 12291
rect 3927 12257 3936 12291
rect 3884 12248 3936 12257
rect 6000 12316 6052 12368
rect 6276 12316 6328 12368
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 9036 12316 9088 12368
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 18420 12427 18472 12436
rect 18420 12393 18429 12427
rect 18429 12393 18463 12427
rect 18463 12393 18472 12427
rect 18420 12384 18472 12393
rect 17408 12316 17460 12368
rect 9772 12248 9824 12300
rect 8116 12180 8168 12232
rect 1676 12155 1728 12164
rect 1676 12121 1685 12155
rect 1685 12121 1719 12155
rect 1719 12121 1728 12155
rect 1676 12112 1728 12121
rect 1952 12112 2004 12164
rect 4252 12112 4304 12164
rect 11060 12155 11112 12164
rect 11060 12121 11069 12155
rect 11069 12121 11103 12155
rect 11103 12121 11112 12155
rect 11060 12112 11112 12121
rect 11520 12180 11572 12232
rect 11428 12112 11480 12164
rect 2964 12044 3016 12096
rect 6276 12044 6328 12096
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 11152 12044 11204 12096
rect 12716 12044 12768 12096
rect 15292 12248 15344 12300
rect 16672 12248 16724 12300
rect 17224 12248 17276 12300
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 14648 12112 14700 12164
rect 15292 12112 15344 12164
rect 14188 12044 14240 12096
rect 16856 12087 16908 12096
rect 16856 12053 16865 12087
rect 16865 12053 16899 12087
rect 16899 12053 16908 12087
rect 16856 12044 16908 12053
rect 17960 12044 18012 12096
rect 3875 11942 3927 11994
rect 3939 11942 3991 11994
rect 4003 11942 4055 11994
rect 4067 11942 4119 11994
rect 4131 11942 4183 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 8534 11942 8586 11994
rect 8598 11942 8650 11994
rect 8662 11942 8714 11994
rect 12937 11942 12989 11994
rect 13001 11942 13053 11994
rect 13065 11942 13117 11994
rect 13129 11942 13181 11994
rect 13193 11942 13245 11994
rect 17468 11942 17520 11994
rect 17532 11942 17584 11994
rect 17596 11942 17648 11994
rect 17660 11942 17712 11994
rect 17724 11942 17776 11994
rect 1676 11840 1728 11892
rect 1952 11883 2004 11892
rect 1952 11849 1961 11883
rect 1961 11849 1995 11883
rect 1995 11849 2004 11883
rect 1952 11840 2004 11849
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 6276 11840 6328 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 9128 11840 9180 11892
rect 9312 11840 9364 11892
rect 9864 11840 9916 11892
rect 11520 11840 11572 11892
rect 13084 11840 13136 11892
rect 13820 11840 13872 11892
rect 15292 11840 15344 11892
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 16856 11840 16908 11892
rect 2044 11704 2096 11756
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2872 11772 2924 11824
rect 3608 11772 3660 11824
rect 2964 11704 3016 11756
rect 3056 11636 3108 11688
rect 4988 11772 5040 11824
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 6184 11704 6236 11756
rect 4252 11636 4304 11688
rect 4436 11679 4488 11688
rect 4436 11645 4445 11679
rect 4445 11645 4479 11679
rect 4479 11645 4488 11679
rect 4436 11636 4488 11645
rect 6920 11772 6972 11824
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 2688 11568 2740 11620
rect 2780 11500 2832 11552
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 12164 11772 12216 11824
rect 16304 11772 16356 11824
rect 9680 11704 9732 11756
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 13360 11704 13412 11756
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 15568 11704 15620 11756
rect 16028 11704 16080 11756
rect 11520 11636 11572 11688
rect 14648 11636 14700 11688
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 9404 11568 9456 11620
rect 10784 11500 10836 11552
rect 12624 11500 12676 11552
rect 12900 11500 12952 11552
rect 3215 11398 3267 11450
rect 3279 11398 3331 11450
rect 3343 11398 3395 11450
rect 3407 11398 3459 11450
rect 3471 11398 3523 11450
rect 7746 11398 7798 11450
rect 7810 11398 7862 11450
rect 7874 11398 7926 11450
rect 7938 11398 7990 11450
rect 8002 11398 8054 11450
rect 12277 11398 12329 11450
rect 12341 11398 12393 11450
rect 12405 11398 12457 11450
rect 12469 11398 12521 11450
rect 12533 11398 12585 11450
rect 16808 11398 16860 11450
rect 16872 11398 16924 11450
rect 16936 11398 16988 11450
rect 17000 11398 17052 11450
rect 17064 11398 17116 11450
rect 3056 11296 3108 11348
rect 6644 11296 6696 11348
rect 9772 11296 9824 11348
rect 12164 11296 12216 11348
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 4436 11092 4488 11144
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 7288 11160 7340 11212
rect 9864 11160 9916 11212
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 11152 11228 11204 11280
rect 12900 11296 12952 11348
rect 13360 11296 13412 11348
rect 12716 11228 12768 11280
rect 11612 11160 11664 11212
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 11152 11092 11204 11144
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 11060 11024 11112 11076
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 14924 11160 14976 11212
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 10416 10999 10468 11008
rect 10416 10965 10425 10999
rect 10425 10965 10459 10999
rect 10459 10965 10468 10999
rect 10416 10956 10468 10965
rect 11244 10956 11296 11008
rect 12716 10956 12768 11008
rect 18880 10999 18932 11008
rect 18880 10965 18889 10999
rect 18889 10965 18923 10999
rect 18923 10965 18932 10999
rect 18880 10956 18932 10965
rect 3875 10854 3927 10906
rect 3939 10854 3991 10906
rect 4003 10854 4055 10906
rect 4067 10854 4119 10906
rect 4131 10854 4183 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 8534 10854 8586 10906
rect 8598 10854 8650 10906
rect 8662 10854 8714 10906
rect 12937 10854 12989 10906
rect 13001 10854 13053 10906
rect 13065 10854 13117 10906
rect 13129 10854 13181 10906
rect 13193 10854 13245 10906
rect 17468 10854 17520 10906
rect 17532 10854 17584 10906
rect 17596 10854 17648 10906
rect 17660 10854 17712 10906
rect 17724 10854 17776 10906
rect 4436 10795 4488 10804
rect 4436 10761 4445 10795
rect 4445 10761 4479 10795
rect 4479 10761 4488 10795
rect 4436 10752 4488 10761
rect 10416 10752 10468 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11152 10752 11204 10804
rect 16212 10752 16264 10804
rect 18328 10752 18380 10804
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 6460 10616 6512 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7472 10616 7524 10668
rect 11060 10616 11112 10668
rect 11336 10659 11388 10668
rect 11336 10625 11337 10659
rect 11337 10625 11371 10659
rect 11371 10625 11388 10659
rect 11336 10616 11388 10625
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 12716 10616 12768 10668
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 17684 10684 17736 10736
rect 16488 10616 16540 10668
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 4252 10548 4304 10600
rect 5080 10548 5132 10600
rect 7656 10548 7708 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 11244 10548 11296 10600
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 13912 10480 13964 10532
rect 16580 10480 16632 10532
rect 3976 10412 4028 10464
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5172 10412 5224 10464
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 14740 10412 14792 10464
rect 17500 10412 17552 10464
rect 3215 10310 3267 10362
rect 3279 10310 3331 10362
rect 3343 10310 3395 10362
rect 3407 10310 3459 10362
rect 3471 10310 3523 10362
rect 7746 10310 7798 10362
rect 7810 10310 7862 10362
rect 7874 10310 7926 10362
rect 7938 10310 7990 10362
rect 8002 10310 8054 10362
rect 12277 10310 12329 10362
rect 12341 10310 12393 10362
rect 12405 10310 12457 10362
rect 12469 10310 12521 10362
rect 12533 10310 12585 10362
rect 16808 10310 16860 10362
rect 16872 10310 16924 10362
rect 16936 10310 16988 10362
rect 17000 10310 17052 10362
rect 17064 10310 17116 10362
rect 3976 10251 4028 10260
rect 3976 10217 3985 10251
rect 3985 10217 4019 10251
rect 4019 10217 4028 10251
rect 3976 10208 4028 10217
rect 4252 10208 4304 10260
rect 4988 10208 5040 10260
rect 7564 10208 7616 10260
rect 4160 10115 4212 10124
rect 4160 10081 4169 10115
rect 4169 10081 4203 10115
rect 4203 10081 4212 10115
rect 4160 10072 4212 10081
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 7288 10072 7340 10124
rect 10600 10208 10652 10260
rect 11704 10208 11756 10260
rect 12624 10208 12676 10260
rect 15292 10208 15344 10260
rect 16028 10140 16080 10192
rect 11152 10072 11204 10124
rect 14280 10072 14332 10124
rect 14740 10072 14792 10124
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 18696 10072 18748 10124
rect 2136 9936 2188 9988
rect 2872 9979 2924 9988
rect 2872 9945 2881 9979
rect 2881 9945 2915 9979
rect 2915 9945 2924 9979
rect 2872 9936 2924 9945
rect 1400 9911 1452 9920
rect 1400 9877 1409 9911
rect 1409 9877 1443 9911
rect 1443 9877 1452 9911
rect 1400 9868 1452 9877
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3608 10004 3660 10056
rect 4528 9936 4580 9988
rect 5172 9936 5224 9988
rect 8300 10004 8352 10056
rect 9036 10004 9088 10056
rect 11244 10004 11296 10056
rect 11704 10004 11756 10056
rect 13636 10004 13688 10056
rect 9220 9936 9272 9988
rect 11612 9936 11664 9988
rect 4804 9868 4856 9920
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 7012 9868 7064 9920
rect 7472 9868 7524 9920
rect 8944 9868 8996 9920
rect 13820 9911 13872 9920
rect 13820 9877 13829 9911
rect 13829 9877 13863 9911
rect 13863 9877 13872 9911
rect 13820 9868 13872 9877
rect 15568 9868 15620 9920
rect 16488 10004 16540 10056
rect 16488 9868 16540 9920
rect 17500 10004 17552 10056
rect 18328 10004 18380 10056
rect 17960 9868 18012 9920
rect 3875 9766 3927 9818
rect 3939 9766 3991 9818
rect 4003 9766 4055 9818
rect 4067 9766 4119 9818
rect 4131 9766 4183 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 8534 9766 8586 9818
rect 8598 9766 8650 9818
rect 8662 9766 8714 9818
rect 12937 9766 12989 9818
rect 13001 9766 13053 9818
rect 13065 9766 13117 9818
rect 13129 9766 13181 9818
rect 13193 9766 13245 9818
rect 17468 9766 17520 9818
rect 17532 9766 17584 9818
rect 17596 9766 17648 9818
rect 17660 9766 17712 9818
rect 17724 9766 17776 9818
rect 2136 9707 2188 9716
rect 2136 9673 2145 9707
rect 2145 9673 2179 9707
rect 2179 9673 2188 9707
rect 2136 9664 2188 9673
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 11152 9664 11204 9716
rect 15660 9664 15712 9716
rect 16488 9664 16540 9716
rect 18696 9664 18748 9716
rect 6000 9596 6052 9648
rect 8944 9596 8996 9648
rect 9404 9639 9456 9648
rect 9404 9605 9413 9639
rect 9413 9605 9447 9639
rect 9447 9605 9456 9639
rect 9404 9596 9456 9605
rect 3240 9528 3292 9580
rect 4712 9528 4764 9580
rect 6828 9528 6880 9580
rect 7656 9528 7708 9580
rect 11244 9528 11296 9580
rect 11888 9596 11940 9648
rect 14096 9596 14148 9648
rect 14280 9596 14332 9648
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 14924 9528 14976 9580
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 2320 9460 2372 9512
rect 5080 9460 5132 9512
rect 6644 9460 6696 9512
rect 2044 9392 2096 9444
rect 4804 9324 4856 9376
rect 5080 9367 5132 9376
rect 5080 9333 5089 9367
rect 5089 9333 5123 9367
rect 5123 9333 5132 9367
rect 5080 9324 5132 9333
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 11520 9460 11572 9512
rect 11704 9460 11756 9512
rect 8300 9392 8352 9444
rect 11152 9392 11204 9444
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 13912 9460 13964 9512
rect 16212 9460 16264 9512
rect 17960 9460 18012 9512
rect 13360 9392 13412 9444
rect 9220 9324 9272 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 11980 9324 12032 9376
rect 13636 9324 13688 9376
rect 3215 9222 3267 9274
rect 3279 9222 3331 9274
rect 3343 9222 3395 9274
rect 3407 9222 3459 9274
rect 3471 9222 3523 9274
rect 7746 9222 7798 9274
rect 7810 9222 7862 9274
rect 7874 9222 7926 9274
rect 7938 9222 7990 9274
rect 8002 9222 8054 9274
rect 12277 9222 12329 9274
rect 12341 9222 12393 9274
rect 12405 9222 12457 9274
rect 12469 9222 12521 9274
rect 12533 9222 12585 9274
rect 16808 9222 16860 9274
rect 16872 9222 16924 9274
rect 16936 9222 16988 9274
rect 17000 9222 17052 9274
rect 17064 9222 17116 9274
rect 7656 9120 7708 9172
rect 11152 9120 11204 9172
rect 11244 9120 11296 9172
rect 12716 9120 12768 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 14096 9120 14148 9172
rect 16212 9120 16264 9172
rect 1400 8984 1452 9036
rect 2412 9027 2464 9036
rect 2412 8993 2421 9027
rect 2421 8993 2455 9027
rect 2455 8993 2464 9027
rect 2412 8984 2464 8993
rect 6644 8984 6696 9036
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2780 8916 2832 8968
rect 4988 8916 5040 8968
rect 9220 8916 9272 8968
rect 9404 8916 9456 8968
rect 10968 8916 11020 8968
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 6460 8848 6512 8900
rect 7012 8848 7064 8900
rect 13544 8916 13596 8968
rect 16580 8984 16632 9036
rect 13820 8916 13872 8968
rect 14924 8916 14976 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 16396 8916 16448 8968
rect 17868 8916 17920 8968
rect 1952 8780 2004 8832
rect 2964 8780 3016 8832
rect 4712 8780 4764 8832
rect 10140 8780 10192 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 3875 8678 3927 8730
rect 3939 8678 3991 8730
rect 4003 8678 4055 8730
rect 4067 8678 4119 8730
rect 4131 8678 4183 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 8534 8678 8586 8730
rect 8598 8678 8650 8730
rect 8662 8678 8714 8730
rect 12937 8678 12989 8730
rect 13001 8678 13053 8730
rect 13065 8678 13117 8730
rect 13129 8678 13181 8730
rect 13193 8678 13245 8730
rect 17468 8678 17520 8730
rect 17532 8678 17584 8730
rect 17596 8678 17648 8730
rect 17660 8678 17712 8730
rect 17724 8678 17776 8730
rect 2412 8576 2464 8628
rect 1952 8372 2004 8424
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 2964 8415 3016 8424
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 3792 8440 3844 8492
rect 5172 8576 5224 8628
rect 6000 8576 6052 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 5540 8508 5592 8560
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 8300 8440 8352 8492
rect 9312 8508 9364 8560
rect 10692 8576 10744 8628
rect 11704 8576 11756 8628
rect 9864 8508 9916 8560
rect 11980 8576 12032 8628
rect 13544 8576 13596 8628
rect 14648 8619 14700 8628
rect 14648 8585 14657 8619
rect 14657 8585 14691 8619
rect 14691 8585 14700 8619
rect 14648 8576 14700 8585
rect 12900 8440 12952 8492
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 12808 8372 12860 8424
rect 13820 8440 13872 8492
rect 14740 8440 14792 8492
rect 18512 8576 18564 8628
rect 15292 8372 15344 8424
rect 15568 8372 15620 8424
rect 16488 8508 16540 8560
rect 17408 8508 17460 8560
rect 16396 8440 16448 8492
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 1768 8279 1820 8288
rect 1768 8245 1777 8279
rect 1777 8245 1811 8279
rect 1811 8245 1820 8279
rect 1768 8236 1820 8245
rect 2872 8236 2924 8288
rect 5080 8236 5132 8288
rect 6000 8279 6052 8288
rect 6000 8245 6009 8279
rect 6009 8245 6043 8279
rect 6043 8245 6052 8279
rect 6000 8236 6052 8245
rect 16580 8304 16632 8356
rect 8760 8236 8812 8288
rect 17592 8236 17644 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 3215 8134 3267 8186
rect 3279 8134 3331 8186
rect 3343 8134 3395 8186
rect 3407 8134 3459 8186
rect 3471 8134 3523 8186
rect 7746 8134 7798 8186
rect 7810 8134 7862 8186
rect 7874 8134 7926 8186
rect 7938 8134 7990 8186
rect 8002 8134 8054 8186
rect 12277 8134 12329 8186
rect 12341 8134 12393 8186
rect 12405 8134 12457 8186
rect 12469 8134 12521 8186
rect 12533 8134 12585 8186
rect 16808 8134 16860 8186
rect 16872 8134 16924 8186
rect 16936 8134 16988 8186
rect 17000 8134 17052 8186
rect 17064 8134 17116 8186
rect 2504 8032 2556 8084
rect 4344 8032 4396 8084
rect 5540 8032 5592 8084
rect 1768 7896 1820 7948
rect 7656 7964 7708 8016
rect 4160 7828 4212 7880
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 7932 7896 7984 7948
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 9864 8032 9916 8084
rect 11520 8032 11572 8084
rect 8760 7896 8812 7948
rect 1400 7760 1452 7812
rect 6644 7760 6696 7812
rect 7012 7803 7064 7812
rect 7012 7769 7021 7803
rect 7021 7769 7055 7803
rect 7055 7769 7064 7803
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 11060 7828 11112 7880
rect 11612 7828 11664 7880
rect 12808 8032 12860 8084
rect 12900 7964 12952 8016
rect 14924 7896 14976 7948
rect 15384 8032 15436 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 17316 8032 17368 8084
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 7012 7760 7064 7769
rect 14004 7828 14056 7880
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 16396 7828 16448 7880
rect 18420 7896 18472 7948
rect 18788 7896 18840 7948
rect 2320 7735 2372 7744
rect 2320 7701 2329 7735
rect 2329 7701 2363 7735
rect 2363 7701 2372 7735
rect 2320 7692 2372 7701
rect 3148 7692 3200 7744
rect 4620 7735 4672 7744
rect 4620 7701 4629 7735
rect 4629 7701 4663 7735
rect 4663 7701 4672 7735
rect 4620 7692 4672 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8208 7692 8260 7744
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 10140 7692 10192 7744
rect 10416 7692 10468 7744
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 14832 7692 14884 7701
rect 15200 7692 15252 7744
rect 17868 7760 17920 7812
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 3875 7590 3927 7642
rect 3939 7590 3991 7642
rect 4003 7590 4055 7642
rect 4067 7590 4119 7642
rect 4131 7590 4183 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 8534 7590 8586 7642
rect 8598 7590 8650 7642
rect 8662 7590 8714 7642
rect 12937 7590 12989 7642
rect 13001 7590 13053 7642
rect 13065 7590 13117 7642
rect 13129 7590 13181 7642
rect 13193 7590 13245 7642
rect 17468 7590 17520 7642
rect 17532 7590 17584 7642
rect 17596 7590 17648 7642
rect 17660 7590 17712 7642
rect 17724 7590 17776 7642
rect 1952 7488 2004 7540
rect 4252 7488 4304 7540
rect 2228 7420 2280 7472
rect 2872 7463 2924 7472
rect 2872 7429 2881 7463
rect 2881 7429 2915 7463
rect 2915 7429 2924 7463
rect 2872 7420 2924 7429
rect 4620 7488 4672 7540
rect 5080 7488 5132 7540
rect 7104 7488 7156 7540
rect 7748 7488 7800 7540
rect 8208 7488 8260 7540
rect 9680 7488 9732 7540
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 10416 7488 10468 7540
rect 14096 7488 14148 7540
rect 14832 7488 14884 7540
rect 14924 7488 14976 7540
rect 17132 7488 17184 7540
rect 18512 7531 18564 7540
rect 18512 7497 18521 7531
rect 18521 7497 18555 7531
rect 18555 7497 18564 7531
rect 18512 7488 18564 7497
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 5540 7352 5592 7404
rect 8944 7420 8996 7472
rect 10324 7463 10376 7472
rect 6000 7284 6052 7336
rect 9404 7284 9456 7336
rect 7932 7216 7984 7268
rect 10324 7429 10333 7463
rect 10333 7429 10367 7463
rect 10367 7429 10376 7463
rect 10324 7420 10376 7429
rect 12900 7420 12952 7472
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 10968 7352 11020 7404
rect 11520 7352 11572 7404
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 15200 7352 15252 7404
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 15384 7284 15436 7336
rect 16580 7284 16632 7336
rect 18788 7352 18840 7404
rect 16672 7148 16724 7200
rect 18604 7148 18656 7200
rect 3215 7046 3267 7098
rect 3279 7046 3331 7098
rect 3343 7046 3395 7098
rect 3407 7046 3459 7098
rect 3471 7046 3523 7098
rect 7746 7046 7798 7098
rect 7810 7046 7862 7098
rect 7874 7046 7926 7098
rect 7938 7046 7990 7098
rect 8002 7046 8054 7098
rect 12277 7046 12329 7098
rect 12341 7046 12393 7098
rect 12405 7046 12457 7098
rect 12469 7046 12521 7098
rect 12533 7046 12585 7098
rect 16808 7046 16860 7098
rect 16872 7046 16924 7098
rect 16936 7046 16988 7098
rect 17000 7046 17052 7098
rect 17064 7046 17116 7098
rect 2228 6944 2280 6996
rect 4252 6944 4304 6996
rect 4988 6944 5040 6996
rect 8944 6944 8996 6996
rect 10600 6944 10652 6996
rect 12900 6987 12952 6996
rect 12900 6953 12909 6987
rect 12909 6953 12943 6987
rect 12943 6953 12952 6987
rect 12900 6944 12952 6953
rect 14004 6944 14056 6996
rect 1860 6808 1912 6860
rect 2596 6808 2648 6860
rect 2688 6672 2740 6724
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 5172 6808 5224 6860
rect 9404 6808 9456 6860
rect 4344 6604 4396 6656
rect 5540 6740 5592 6792
rect 10416 6740 10468 6792
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 15200 6876 15252 6928
rect 15292 6876 15344 6928
rect 13728 6808 13780 6860
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 14096 6740 14148 6792
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 15476 6740 15528 6792
rect 15568 6783 15620 6792
rect 15568 6749 15577 6783
rect 15577 6749 15611 6783
rect 15611 6749 15620 6783
rect 15568 6740 15620 6749
rect 15936 6672 15988 6724
rect 5448 6604 5500 6656
rect 8760 6604 8812 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 11796 6604 11848 6656
rect 12624 6604 12676 6656
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 15568 6604 15620 6656
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 16028 6604 16080 6656
rect 16856 6808 16908 6860
rect 16764 6740 16816 6792
rect 16580 6604 16632 6656
rect 17040 6604 17092 6656
rect 3875 6502 3927 6554
rect 3939 6502 3991 6554
rect 4003 6502 4055 6554
rect 4067 6502 4119 6554
rect 4131 6502 4183 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 8534 6502 8586 6554
rect 8598 6502 8650 6554
rect 8662 6502 8714 6554
rect 12937 6502 12989 6554
rect 13001 6502 13053 6554
rect 13065 6502 13117 6554
rect 13129 6502 13181 6554
rect 13193 6502 13245 6554
rect 17468 6502 17520 6554
rect 17532 6502 17584 6554
rect 17596 6502 17648 6554
rect 17660 6502 17712 6554
rect 17724 6502 17776 6554
rect 3056 6400 3108 6452
rect 3148 6400 3200 6452
rect 2228 6332 2280 6384
rect 5172 6400 5224 6452
rect 9680 6400 9732 6452
rect 14648 6400 14700 6452
rect 7656 6332 7708 6384
rect 9496 6332 9548 6384
rect 3792 6196 3844 6248
rect 7012 6264 7064 6316
rect 12808 6332 12860 6384
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 2136 6060 2188 6112
rect 5264 6196 5316 6248
rect 9312 6196 9364 6248
rect 11612 6264 11664 6316
rect 15568 6332 15620 6384
rect 16764 6332 16816 6384
rect 17040 6332 17092 6384
rect 15844 6264 15896 6316
rect 16304 6264 16356 6316
rect 18788 6400 18840 6452
rect 17408 6375 17460 6384
rect 17408 6341 17417 6375
rect 17417 6341 17451 6375
rect 17451 6341 17460 6375
rect 17408 6332 17460 6341
rect 18420 6332 18472 6384
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 18144 6196 18196 6248
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 9220 6060 9272 6112
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10692 6060 10744 6069
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 16212 6128 16264 6180
rect 16856 6128 16908 6180
rect 15936 6060 15988 6112
rect 17868 6060 17920 6112
rect 3215 5958 3267 6010
rect 3279 5958 3331 6010
rect 3343 5958 3395 6010
rect 3407 5958 3459 6010
rect 3471 5958 3523 6010
rect 7746 5958 7798 6010
rect 7810 5958 7862 6010
rect 7874 5958 7926 6010
rect 7938 5958 7990 6010
rect 8002 5958 8054 6010
rect 12277 5958 12329 6010
rect 12341 5958 12393 6010
rect 12405 5958 12457 6010
rect 12469 5958 12521 6010
rect 12533 5958 12585 6010
rect 16808 5958 16860 6010
rect 16872 5958 16924 6010
rect 16936 5958 16988 6010
rect 17000 5958 17052 6010
rect 17064 5958 17116 6010
rect 1400 5856 1452 5908
rect 2228 5856 2280 5908
rect 2596 5720 2648 5772
rect 4252 5720 4304 5772
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 2504 5559 2556 5568
rect 2504 5525 2513 5559
rect 2513 5525 2547 5559
rect 2547 5525 2556 5559
rect 2504 5516 2556 5525
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 4620 5652 4672 5704
rect 3792 5584 3844 5636
rect 5172 5695 5224 5704
rect 5172 5661 5181 5695
rect 5181 5661 5215 5695
rect 5215 5661 5224 5695
rect 5172 5652 5224 5661
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 9220 5856 9272 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 11520 5856 11572 5908
rect 12808 5856 12860 5908
rect 16672 5856 16724 5908
rect 17408 5856 17460 5908
rect 18420 5856 18472 5908
rect 8760 5788 8812 5840
rect 2688 5516 2740 5568
rect 4896 5559 4948 5568
rect 4896 5525 4905 5559
rect 4905 5525 4939 5559
rect 4939 5525 4948 5559
rect 4896 5516 4948 5525
rect 5356 5584 5408 5636
rect 6920 5584 6972 5636
rect 9220 5652 9272 5704
rect 11888 5788 11940 5840
rect 10968 5720 11020 5772
rect 11704 5720 11756 5772
rect 16028 5788 16080 5840
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 12624 5652 12676 5704
rect 10692 5584 10744 5636
rect 16212 5695 16264 5704
rect 16212 5661 16228 5695
rect 16228 5661 16262 5695
rect 16262 5661 16264 5695
rect 16212 5652 16264 5661
rect 17868 5652 17920 5704
rect 11980 5516 12032 5568
rect 12624 5516 12676 5568
rect 3875 5414 3927 5466
rect 3939 5414 3991 5466
rect 4003 5414 4055 5466
rect 4067 5414 4119 5466
rect 4131 5414 4183 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 8534 5414 8586 5466
rect 8598 5414 8650 5466
rect 8662 5414 8714 5466
rect 12937 5414 12989 5466
rect 13001 5414 13053 5466
rect 13065 5414 13117 5466
rect 13129 5414 13181 5466
rect 13193 5414 13245 5466
rect 17468 5414 17520 5466
rect 17532 5414 17584 5466
rect 17596 5414 17648 5466
rect 17660 5414 17712 5466
rect 17724 5414 17776 5466
rect 2964 5312 3016 5364
rect 4896 5312 4948 5364
rect 6920 5312 6972 5364
rect 5724 5244 5776 5296
rect 9588 5312 9640 5364
rect 11612 5312 11664 5364
rect 14096 5312 14148 5364
rect 14648 5312 14700 5364
rect 16304 5312 16356 5364
rect 4160 5151 4212 5160
rect 4160 5117 4169 5151
rect 4169 5117 4203 5151
rect 4203 5117 4212 5151
rect 4160 5108 4212 5117
rect 4252 5108 4304 5160
rect 1768 5040 1820 5092
rect 2320 5040 2372 5092
rect 5356 5108 5408 5160
rect 5448 5108 5500 5160
rect 7012 5176 7064 5228
rect 9680 5244 9732 5296
rect 8760 5108 8812 5160
rect 10968 5176 11020 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 12624 5244 12676 5296
rect 13268 5244 13320 5296
rect 15108 5244 15160 5296
rect 9312 5108 9364 5160
rect 11704 5108 11756 5160
rect 11980 5151 12032 5160
rect 11980 5117 11989 5151
rect 11989 5117 12023 5151
rect 12023 5117 12032 5151
rect 11980 5108 12032 5117
rect 14924 5108 14976 5160
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 3215 4870 3267 4922
rect 3279 4870 3331 4922
rect 3343 4870 3395 4922
rect 3407 4870 3459 4922
rect 3471 4870 3523 4922
rect 7746 4870 7798 4922
rect 7810 4870 7862 4922
rect 7874 4870 7926 4922
rect 7938 4870 7990 4922
rect 8002 4870 8054 4922
rect 12277 4870 12329 4922
rect 12341 4870 12393 4922
rect 12405 4870 12457 4922
rect 12469 4870 12521 4922
rect 12533 4870 12585 4922
rect 16808 4870 16860 4922
rect 16872 4870 16924 4922
rect 16936 4870 16988 4922
rect 17000 4870 17052 4922
rect 17064 4870 17116 4922
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 4160 4768 4212 4820
rect 5724 4811 5776 4820
rect 5724 4777 5733 4811
rect 5733 4777 5767 4811
rect 5767 4777 5776 4811
rect 5724 4768 5776 4777
rect 6184 4768 6236 4820
rect 9680 4768 9732 4820
rect 13268 4768 13320 4820
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 2504 4632 2556 4684
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 5448 4564 5500 4616
rect 8760 4564 8812 4616
rect 12716 4564 12768 4616
rect 14924 4564 14976 4616
rect 2780 4496 2832 4548
rect 3875 4326 3927 4378
rect 3939 4326 3991 4378
rect 4003 4326 4055 4378
rect 4067 4326 4119 4378
rect 4131 4326 4183 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 8534 4326 8586 4378
rect 8598 4326 8650 4378
rect 8662 4326 8714 4378
rect 12937 4326 12989 4378
rect 13001 4326 13053 4378
rect 13065 4326 13117 4378
rect 13129 4326 13181 4378
rect 13193 4326 13245 4378
rect 17468 4326 17520 4378
rect 17532 4326 17584 4378
rect 17596 4326 17648 4378
rect 17660 4326 17712 4378
rect 17724 4326 17776 4378
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 14924 4224 14976 4276
rect 15292 4199 15344 4208
rect 15292 4165 15301 4199
rect 15301 4165 15335 4199
rect 15335 4165 15344 4199
rect 15292 4156 15344 4165
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 3215 3782 3267 3834
rect 3279 3782 3331 3834
rect 3343 3782 3395 3834
rect 3407 3782 3459 3834
rect 3471 3782 3523 3834
rect 7746 3782 7798 3834
rect 7810 3782 7862 3834
rect 7874 3782 7926 3834
rect 7938 3782 7990 3834
rect 8002 3782 8054 3834
rect 12277 3782 12329 3834
rect 12341 3782 12393 3834
rect 12405 3782 12457 3834
rect 12469 3782 12521 3834
rect 12533 3782 12585 3834
rect 16808 3782 16860 3834
rect 16872 3782 16924 3834
rect 16936 3782 16988 3834
rect 17000 3782 17052 3834
rect 17064 3782 17116 3834
rect 3875 3238 3927 3290
rect 3939 3238 3991 3290
rect 4003 3238 4055 3290
rect 4067 3238 4119 3290
rect 4131 3238 4183 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 8534 3238 8586 3290
rect 8598 3238 8650 3290
rect 8662 3238 8714 3290
rect 12937 3238 12989 3290
rect 13001 3238 13053 3290
rect 13065 3238 13117 3290
rect 13129 3238 13181 3290
rect 13193 3238 13245 3290
rect 17468 3238 17520 3290
rect 17532 3238 17584 3290
rect 17596 3238 17648 3290
rect 17660 3238 17712 3290
rect 17724 3238 17776 3290
rect 3215 2694 3267 2746
rect 3279 2694 3331 2746
rect 3343 2694 3395 2746
rect 3407 2694 3459 2746
rect 3471 2694 3523 2746
rect 7746 2694 7798 2746
rect 7810 2694 7862 2746
rect 7874 2694 7926 2746
rect 7938 2694 7990 2746
rect 8002 2694 8054 2746
rect 12277 2694 12329 2746
rect 12341 2694 12393 2746
rect 12405 2694 12457 2746
rect 12469 2694 12521 2746
rect 12533 2694 12585 2746
rect 16808 2694 16860 2746
rect 16872 2694 16924 2746
rect 16936 2694 16988 2746
rect 17000 2694 17052 2746
rect 17064 2694 17116 2746
rect 15292 2592 15344 2644
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 3875 2150 3927 2202
rect 3939 2150 3991 2202
rect 4003 2150 4055 2202
rect 4067 2150 4119 2202
rect 4131 2150 4183 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 8534 2150 8586 2202
rect 8598 2150 8650 2202
rect 8662 2150 8714 2202
rect 12937 2150 12989 2202
rect 13001 2150 13053 2202
rect 13065 2150 13117 2202
rect 13129 2150 13181 2202
rect 13193 2150 13245 2202
rect 17468 2150 17520 2202
rect 17532 2150 17584 2202
rect 17596 2150 17648 2202
rect 17660 2150 17712 2202
rect 17724 2150 17776 2202
<< metal2 >>
rect 1582 21714 1638 22514
rect 2134 21714 2190 22514
rect 2686 21714 2742 22514
rect 3238 21714 3294 22514
rect 3790 21714 3846 22514
rect 4342 21714 4398 22514
rect 4894 21714 4950 22514
rect 5446 21714 5502 22514
rect 5998 21714 6054 22514
rect 6550 21714 6606 22514
rect 7102 21714 7158 22514
rect 7654 21714 7710 22514
rect 8206 21714 8262 22514
rect 8758 21714 8814 22514
rect 9310 21714 9366 22514
rect 9862 21714 9918 22514
rect 10414 21714 10470 22514
rect 10966 21714 11022 22514
rect 11518 21714 11574 22514
rect 12070 21714 12126 22514
rect 12622 21714 12678 22514
rect 13174 21714 13230 22514
rect 13726 21714 13782 22514
rect 14278 21714 14334 22514
rect 14830 21842 14886 22514
rect 14830 21814 15148 21842
rect 14830 21714 14886 21814
rect 1596 19854 1624 21714
rect 2148 19854 2176 21714
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 2136 19848 2188 19854
rect 2700 19836 2728 21714
rect 3252 20346 3280 21714
rect 3068 20318 3280 20346
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 2780 19848 2832 19854
rect 2700 19808 2780 19836
rect 2136 19790 2188 19796
rect 2780 19790 2832 19796
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1780 18290 1808 18566
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 16697 980 17138
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 938 16688 994 16697
rect 938 16623 994 16632
rect 1596 16182 1624 16934
rect 1584 16176 1636 16182
rect 1584 16118 1636 16124
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1412 12306 1440 14894
rect 1688 14618 1716 14894
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 11898 1716 12106
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9042 1440 9862
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 7818 1440 8978
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1780 7954 1808 8230
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1400 7812 1452 7818
rect 1400 7754 1452 7760
rect 1872 6866 1900 19654
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 14414 2084 17138
rect 2148 15722 2176 19654
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2792 19258 2820 19314
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2700 19230 2820 19258
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2608 18698 2636 19178
rect 2700 18970 2728 19230
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2700 17338 2728 18906
rect 2792 18630 2820 19110
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2884 18222 2912 19246
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2884 17678 2912 18158
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2976 17490 3004 19926
rect 3068 19854 3096 20318
rect 3215 20156 3523 20165
rect 3215 20154 3221 20156
rect 3277 20154 3301 20156
rect 3357 20154 3381 20156
rect 3437 20154 3461 20156
rect 3517 20154 3523 20156
rect 3277 20102 3279 20154
rect 3459 20102 3461 20154
rect 3215 20100 3221 20102
rect 3277 20100 3301 20102
rect 3357 20100 3381 20102
rect 3437 20100 3461 20102
rect 3517 20100 3523 20102
rect 3215 20091 3523 20100
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3160 19394 3188 19994
rect 3804 19854 3832 21714
rect 4356 19854 4384 21714
rect 4908 19854 4936 21714
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4896 19848 4948 19854
rect 5460 19836 5488 21714
rect 6012 19854 6040 21714
rect 6564 20058 6592 21714
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 7116 19854 7144 21714
rect 7668 19854 7696 21714
rect 7746 20156 8054 20165
rect 7746 20154 7752 20156
rect 7808 20154 7832 20156
rect 7888 20154 7912 20156
rect 7968 20154 7992 20156
rect 8048 20154 8054 20156
rect 7808 20102 7810 20154
rect 7990 20102 7992 20154
rect 7746 20100 7752 20102
rect 7808 20100 7832 20102
rect 7888 20100 7912 20102
rect 7968 20100 7992 20102
rect 8048 20100 8054 20102
rect 7746 20091 8054 20100
rect 5540 19848 5592 19854
rect 5460 19808 5540 19836
rect 4896 19790 4948 19796
rect 5540 19790 5592 19796
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7656 19848 7708 19854
rect 8220 19836 8248 21714
rect 8772 19854 8800 21714
rect 9220 19984 9272 19990
rect 9220 19926 9272 19932
rect 8300 19848 8352 19854
rect 8220 19808 8300 19836
rect 7656 19790 7708 19796
rect 8300 19790 8352 19796
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 3068 19366 3188 19394
rect 3068 19310 3096 19366
rect 3528 19334 3556 19654
rect 3875 19612 4183 19621
rect 3875 19610 3881 19612
rect 3937 19610 3961 19612
rect 4017 19610 4041 19612
rect 4097 19610 4121 19612
rect 4177 19610 4183 19612
rect 3937 19558 3939 19610
rect 4119 19558 4121 19610
rect 3875 19556 3881 19558
rect 3937 19556 3961 19558
rect 4017 19556 4041 19558
rect 4097 19556 4121 19558
rect 4177 19556 4183 19558
rect 3875 19547 4183 19556
rect 3884 19372 3936 19378
rect 3056 19304 3108 19310
rect 3528 19306 3740 19334
rect 3884 19314 3936 19320
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 3056 19246 3108 19252
rect 3068 17762 3096 19246
rect 3215 19068 3523 19077
rect 3215 19066 3221 19068
rect 3277 19066 3301 19068
rect 3357 19066 3381 19068
rect 3437 19066 3461 19068
rect 3517 19066 3523 19068
rect 3277 19014 3279 19066
rect 3459 19014 3461 19066
rect 3215 19012 3221 19014
rect 3277 19012 3301 19014
rect 3357 19012 3381 19014
rect 3437 19012 3461 19014
rect 3517 19012 3523 19014
rect 3215 19003 3523 19012
rect 3712 18986 3740 19306
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3620 18958 3740 18986
rect 3620 18952 3648 18958
rect 3528 18924 3648 18952
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3160 18290 3188 18702
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3528 18068 3556 18924
rect 3700 18896 3752 18902
rect 3700 18838 3752 18844
rect 3712 18290 3740 18838
rect 3804 18426 3832 19110
rect 3896 18698 3924 19314
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18970 4016 19246
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3884 18692 3936 18698
rect 3884 18634 3936 18640
rect 3875 18524 4183 18533
rect 3875 18522 3881 18524
rect 3937 18522 3961 18524
rect 4017 18522 4041 18524
rect 4097 18522 4121 18524
rect 4177 18522 4183 18524
rect 3937 18470 3939 18522
rect 4119 18470 4121 18522
rect 3875 18468 3881 18470
rect 3937 18468 3961 18470
rect 4017 18468 4041 18470
rect 4097 18468 4121 18470
rect 4177 18468 4183 18470
rect 3875 18459 4183 18468
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 4264 18358 4292 19314
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4356 18426 4384 19246
rect 4436 19236 4488 19242
rect 4436 19178 4488 19184
rect 4448 18902 4476 19178
rect 4436 18896 4488 18902
rect 4436 18838 4488 18844
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4252 18352 4304 18358
rect 4252 18294 4304 18300
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 3528 18040 3648 18068
rect 3215 17980 3523 17989
rect 3215 17978 3221 17980
rect 3277 17978 3301 17980
rect 3357 17978 3381 17980
rect 3437 17978 3461 17980
rect 3517 17978 3523 17980
rect 3277 17926 3279 17978
rect 3459 17926 3461 17978
rect 3215 17924 3221 17926
rect 3277 17924 3301 17926
rect 3357 17924 3381 17926
rect 3437 17924 3461 17926
rect 3517 17924 3523 17926
rect 3215 17915 3523 17924
rect 3068 17734 3188 17762
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2792 17462 3004 17490
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 16522 2268 16934
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2148 15694 2360 15722
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2148 14550 2176 15030
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2240 14482 2268 15506
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 13326 2084 14350
rect 2240 13870 2268 14418
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2332 13682 2360 15694
rect 2700 14414 2728 17070
rect 2792 16538 2820 17462
rect 3068 17134 3096 17614
rect 3160 17338 3188 17734
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16658 2912 16934
rect 3215 16892 3523 16901
rect 3215 16890 3221 16892
rect 3277 16890 3301 16892
rect 3357 16890 3381 16892
rect 3437 16890 3461 16892
rect 3517 16890 3523 16892
rect 3277 16838 3279 16890
rect 3459 16838 3461 16890
rect 3215 16836 3221 16838
rect 3277 16836 3301 16838
rect 3357 16836 3381 16838
rect 3437 16836 3461 16838
rect 3517 16836 3523 16838
rect 3215 16827 3523 16836
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2792 16510 2912 16538
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 15570 2820 16390
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2792 14482 2820 14826
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2688 14408 2740 14414
rect 2740 14356 2820 14362
rect 2688 14350 2820 14356
rect 2700 14334 2820 14350
rect 2240 13654 2360 13682
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1964 11898 1992 12106
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2056 11762 2084 13262
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 9450 2084 11698
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2148 9722 2176 9930
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 2240 9330 2268 13654
rect 2686 12880 2742 12889
rect 2686 12815 2688 12824
rect 2740 12815 2742 12824
rect 2688 12786 2740 12792
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2332 11370 2360 11698
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2700 11370 2728 11562
rect 2792 11558 2820 14334
rect 2884 11830 2912 16510
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3068 14482 3096 16390
rect 3215 15804 3523 15813
rect 3215 15802 3221 15804
rect 3277 15802 3301 15804
rect 3357 15802 3381 15804
rect 3437 15802 3461 15804
rect 3517 15802 3523 15804
rect 3277 15750 3279 15802
rect 3459 15750 3461 15802
rect 3215 15748 3221 15750
rect 3277 15748 3301 15750
rect 3357 15748 3381 15750
rect 3437 15748 3461 15750
rect 3517 15748 3523 15750
rect 3215 15739 3523 15748
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3160 15162 3188 15438
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3436 15026 3464 15506
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3215 14716 3523 14725
rect 3215 14714 3221 14716
rect 3277 14714 3301 14716
rect 3357 14714 3381 14716
rect 3437 14714 3461 14716
rect 3517 14714 3523 14716
rect 3277 14662 3279 14714
rect 3459 14662 3461 14714
rect 3215 14660 3221 14662
rect 3277 14660 3301 14662
rect 3357 14660 3381 14662
rect 3437 14660 3461 14662
rect 3517 14660 3523 14662
rect 3215 14651 3523 14660
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 14074 3096 14214
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3215 13628 3523 13637
rect 3215 13626 3221 13628
rect 3277 13626 3301 13628
rect 3357 13626 3381 13628
rect 3437 13626 3461 13628
rect 3517 13626 3523 13628
rect 3277 13574 3279 13626
rect 3459 13574 3461 13626
rect 3215 13572 3221 13574
rect 3277 13572 3301 13574
rect 3357 13572 3381 13574
rect 3437 13572 3461 13574
rect 3517 13572 3523 13574
rect 3215 13563 3523 13572
rect 3620 12866 3648 18040
rect 3804 17678 3832 18226
rect 4448 18222 4476 18702
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3804 16590 3832 17614
rect 3875 17436 4183 17445
rect 3875 17434 3881 17436
rect 3937 17434 3961 17436
rect 4017 17434 4041 17436
rect 4097 17434 4121 17436
rect 4177 17434 4183 17436
rect 3937 17382 3939 17434
rect 4119 17382 4121 17434
rect 3875 17380 3881 17382
rect 3937 17380 3961 17382
rect 4017 17380 4041 17382
rect 4097 17380 4121 17382
rect 4177 17380 4183 17382
rect 3875 17371 4183 17380
rect 4540 16674 4568 19654
rect 4632 17218 4660 19654
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4724 18970 4752 19246
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4908 18766 4936 19110
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4816 17338 4844 18022
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4632 17190 4844 17218
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4356 16646 4568 16674
rect 4632 16658 4660 16934
rect 4620 16652 4672 16658
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3875 16348 4183 16357
rect 3875 16346 3881 16348
rect 3937 16346 3961 16348
rect 4017 16346 4041 16348
rect 4097 16346 4121 16348
rect 4177 16346 4183 16348
rect 3937 16294 3939 16346
rect 4119 16294 4121 16346
rect 3875 16292 3881 16294
rect 3937 16292 3961 16294
rect 4017 16292 4041 16294
rect 4097 16292 4121 16294
rect 4177 16292 4183 16294
rect 3875 16283 4183 16292
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15026 3832 15302
rect 3875 15260 4183 15269
rect 3875 15258 3881 15260
rect 3937 15258 3961 15260
rect 4017 15258 4041 15260
rect 4097 15258 4121 15260
rect 4177 15258 4183 15260
rect 3937 15206 3939 15258
rect 4119 15206 4121 15258
rect 3875 15204 3881 15206
rect 3937 15204 3961 15206
rect 4017 15204 4041 15206
rect 4097 15204 4121 15206
rect 4177 15204 4183 15206
rect 3875 15195 4183 15204
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3712 13802 3740 14282
rect 3700 13796 3752 13802
rect 3700 13738 3752 13744
rect 3804 12968 3832 14350
rect 3875 14172 4183 14181
rect 3875 14170 3881 14172
rect 3937 14170 3961 14172
rect 4017 14170 4041 14172
rect 4097 14170 4121 14172
rect 4177 14170 4183 14172
rect 3937 14118 3939 14170
rect 4119 14118 4121 14170
rect 3875 14116 3881 14118
rect 3937 14116 3961 14118
rect 4017 14116 4041 14118
rect 4097 14116 4121 14118
rect 4177 14116 4183 14118
rect 3875 14107 4183 14116
rect 4264 14006 4292 15846
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 3875 13084 4183 13093
rect 3875 13082 3881 13084
rect 3937 13082 3961 13084
rect 4017 13082 4041 13084
rect 4097 13082 4121 13084
rect 4177 13082 4183 13084
rect 3937 13030 3939 13082
rect 4119 13030 4121 13082
rect 3875 13028 3881 13030
rect 3937 13028 3961 13030
rect 4017 13028 4041 13030
rect 4097 13028 4121 13030
rect 4177 13028 4183 13030
rect 3875 13019 4183 13028
rect 3804 12940 3924 12968
rect 3620 12838 3832 12866
rect 3215 12540 3523 12549
rect 3215 12538 3221 12540
rect 3277 12538 3301 12540
rect 3357 12538 3381 12540
rect 3437 12538 3461 12540
rect 3517 12538 3523 12540
rect 3277 12486 3279 12538
rect 3459 12486 3461 12538
rect 3215 12484 3221 12486
rect 3277 12484 3301 12486
rect 3357 12484 3381 12486
rect 3437 12484 3461 12486
rect 3517 12484 3523 12486
rect 3215 12475 3523 12484
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2976 11762 3004 12038
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2332 11342 2728 11370
rect 2332 9518 2360 11342
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2148 9302 2268 9330
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8430 1992 8774
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 7546 1992 8366
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2148 6118 2176 9302
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 8634 2452 8978
rect 2792 8974 2820 11494
rect 2976 11218 3004 11698
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3068 11354 3096 11630
rect 3215 11452 3523 11461
rect 3215 11450 3221 11452
rect 3277 11450 3301 11452
rect 3357 11450 3381 11452
rect 3437 11450 3461 11452
rect 3517 11450 3523 11452
rect 3277 11398 3279 11450
rect 3459 11398 3461 11450
rect 3215 11396 3221 11398
rect 3277 11396 3301 11398
rect 3357 11396 3381 11398
rect 3437 11396 3461 11398
rect 3517 11396 3523 11398
rect 3215 11387 3523 11396
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3215 10364 3523 10373
rect 3215 10362 3221 10364
rect 3277 10362 3301 10364
rect 3357 10362 3381 10364
rect 3437 10362 3461 10364
rect 3517 10362 3523 10364
rect 3277 10310 3279 10362
rect 3459 10310 3461 10362
rect 3215 10308 3221 10310
rect 3277 10308 3301 10310
rect 3357 10308 3381 10310
rect 3437 10308 3461 10310
rect 3517 10308 3523 10310
rect 3215 10299 3523 10308
rect 3620 10062 3648 11766
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2884 9722 2912 9930
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3252 9586 3280 9862
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3215 9276 3523 9285
rect 3215 9274 3221 9276
rect 3277 9274 3301 9276
rect 3357 9274 3381 9276
rect 3437 9274 3461 9276
rect 3517 9274 3523 9276
rect 3277 9222 3279 9274
rect 3459 9222 3461 9274
rect 3215 9220 3221 9222
rect 3277 9220 3301 9222
rect 3357 9220 3381 9222
rect 3437 9220 3461 9222
rect 3517 9220 3523 9222
rect 3215 9211 3523 9220
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2516 8090 2544 8910
rect 2792 8412 2820 8910
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8430 3004 8774
rect 3804 8498 3832 12838
rect 3896 12646 3924 12940
rect 4264 12918 4292 13670
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3896 12306 3924 12582
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 3875 11996 4183 12005
rect 3875 11994 3881 11996
rect 3937 11994 3961 11996
rect 4017 11994 4041 11996
rect 4097 11994 4121 11996
rect 4177 11994 4183 11996
rect 3937 11942 3939 11994
rect 4119 11942 4121 11994
rect 3875 11940 3881 11942
rect 3937 11940 3961 11942
rect 4017 11940 4041 11942
rect 4097 11940 4121 11942
rect 4177 11940 4183 11942
rect 3875 11931 4183 11940
rect 4264 11898 4292 12106
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 3875 10908 4183 10917
rect 3875 10906 3881 10908
rect 3937 10906 3961 10908
rect 4017 10906 4041 10908
rect 4097 10906 4121 10908
rect 4177 10906 4183 10908
rect 3937 10854 3939 10906
rect 4119 10854 4121 10906
rect 3875 10852 3881 10854
rect 3937 10852 3961 10854
rect 4017 10852 4041 10854
rect 4097 10852 4121 10854
rect 4177 10852 4183 10854
rect 3875 10843 4183 10852
rect 4264 10606 4292 11630
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 3988 10266 4016 10406
rect 4264 10266 4292 10406
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4172 10010 4200 10066
rect 4172 9982 4292 10010
rect 3875 9820 4183 9829
rect 3875 9818 3881 9820
rect 3937 9818 3961 9820
rect 4017 9818 4041 9820
rect 4097 9818 4121 9820
rect 4177 9818 4183 9820
rect 3937 9766 3939 9818
rect 4119 9766 4121 9818
rect 3875 9764 3881 9766
rect 3937 9764 3961 9766
rect 4017 9764 4041 9766
rect 4097 9764 4121 9766
rect 4177 9764 4183 9766
rect 3875 9755 4183 9764
rect 3875 8732 4183 8741
rect 3875 8730 3881 8732
rect 3937 8730 3961 8732
rect 4017 8730 4041 8732
rect 4097 8730 4121 8732
rect 4177 8730 4183 8732
rect 3937 8678 3939 8730
rect 4119 8678 4121 8730
rect 3875 8676 3881 8678
rect 3937 8676 3961 8678
rect 4017 8676 4041 8678
rect 4097 8676 4121 8678
rect 4177 8676 4183 8678
rect 3875 8667 4183 8676
rect 4264 8498 4292 9982
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 2872 8424 2924 8430
rect 2792 8384 2872 8412
rect 2872 8366 2924 8372
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 4158 8256 4214 8265
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2240 7002 2268 7414
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 1412 5914 1440 6054
rect 2240 5914 2268 6326
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 2332 5098 2360 7686
rect 2884 7478 2912 8230
rect 3215 8188 3523 8197
rect 4158 8191 4214 8200
rect 3215 8186 3221 8188
rect 3277 8186 3301 8188
rect 3357 8186 3381 8188
rect 3437 8186 3461 8188
rect 3517 8186 3523 8188
rect 3277 8134 3279 8186
rect 3459 8134 3461 8186
rect 3215 8132 3221 8134
rect 3277 8132 3301 8134
rect 3357 8132 3381 8134
rect 3437 8132 3461 8134
rect 3517 8132 3523 8134
rect 3215 8123 3523 8132
rect 4172 7886 4200 8191
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 3160 7410 3188 7686
rect 3875 7644 4183 7653
rect 3875 7642 3881 7644
rect 3937 7642 3961 7644
rect 4017 7642 4041 7644
rect 4097 7642 4121 7644
rect 4177 7642 4183 7644
rect 3937 7590 3939 7642
rect 4119 7590 4121 7642
rect 3875 7588 3881 7590
rect 3937 7588 3961 7590
rect 4017 7588 4041 7590
rect 4097 7588 4121 7590
rect 4177 7588 4183 7590
rect 3875 7579 4183 7588
rect 4264 7546 4292 8434
rect 4356 8090 4384 16646
rect 4620 16594 4672 16600
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4540 16250 4568 16458
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12866 4660 13330
rect 4448 12838 4660 12866
rect 4448 11694 4476 12838
rect 4816 12730 4844 17190
rect 4908 16998 4936 18702
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 5000 14278 5028 19654
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5368 18222 5396 18770
rect 5552 18426 5580 18838
rect 5828 18426 5856 19314
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6196 18834 6224 19110
rect 6380 18902 6408 19654
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 6012 18290 6040 18634
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5092 16998 5120 17206
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 15910 5120 16934
rect 5276 16182 5304 17070
rect 5736 17066 5764 17546
rect 5920 17202 5948 18022
rect 6460 17604 6512 17610
rect 6460 17546 6512 17552
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5920 16998 5948 17138
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 6472 16794 6500 17546
rect 6564 17338 6592 19654
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18426 6684 18770
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 5552 16250 5580 16390
rect 6288 16250 6316 16390
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5552 14618 5580 16050
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 6288 14346 6316 15302
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4908 13274 4936 13942
rect 6288 13870 6316 14282
rect 6380 13870 6408 16050
rect 6472 15978 6500 16390
rect 6840 16182 6868 19314
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 16998 6960 18226
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6472 15502 6500 15914
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6932 15434 6960 16934
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6932 15026 6960 15370
rect 7208 15162 7236 19654
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7300 18970 7328 19246
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7392 16538 7420 19654
rect 8406 19612 8714 19621
rect 8406 19610 8412 19612
rect 8468 19610 8492 19612
rect 8548 19610 8572 19612
rect 8628 19610 8652 19612
rect 8708 19610 8714 19612
rect 8468 19558 8470 19610
rect 8650 19558 8652 19610
rect 8406 19556 8412 19558
rect 8468 19556 8492 19558
rect 8548 19556 8572 19558
rect 8628 19556 8652 19558
rect 8708 19556 8714 19558
rect 8406 19547 8714 19556
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 7746 19068 8054 19077
rect 7746 19066 7752 19068
rect 7808 19066 7832 19068
rect 7888 19066 7912 19068
rect 7968 19066 7992 19068
rect 8048 19066 8054 19068
rect 7808 19014 7810 19066
rect 7990 19014 7992 19066
rect 7746 19012 7752 19014
rect 7808 19012 7832 19014
rect 7888 19012 7912 19014
rect 7968 19012 7992 19014
rect 8048 19012 8054 19014
rect 7746 19003 8054 19012
rect 8864 18970 8892 19110
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 7576 18222 7604 18702
rect 8496 18630 8524 18702
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8406 18524 8714 18533
rect 8406 18522 8412 18524
rect 8468 18522 8492 18524
rect 8548 18522 8572 18524
rect 8628 18522 8652 18524
rect 8708 18522 8714 18524
rect 8468 18470 8470 18522
rect 8650 18470 8652 18522
rect 8406 18468 8412 18470
rect 8468 18468 8492 18470
rect 8548 18468 8572 18470
rect 8628 18468 8652 18470
rect 8708 18468 8714 18470
rect 8406 18459 8714 18468
rect 8864 18290 8892 18906
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7576 17882 7604 18158
rect 7746 17980 8054 17989
rect 7746 17978 7752 17980
rect 7808 17978 7832 17980
rect 7888 17978 7912 17980
rect 7968 17978 7992 17980
rect 8048 17978 8054 17980
rect 7808 17926 7810 17978
rect 7990 17926 7992 17978
rect 7746 17924 7752 17926
rect 7808 17924 7832 17926
rect 7888 17924 7912 17926
rect 7968 17924 7992 17926
rect 8048 17924 8054 17926
rect 7746 17915 8054 17924
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 8406 17436 8714 17445
rect 8406 17434 8412 17436
rect 8468 17434 8492 17436
rect 8548 17434 8572 17436
rect 8628 17434 8652 17436
rect 8708 17434 8714 17436
rect 8468 17382 8470 17434
rect 8650 17382 8652 17434
rect 8406 17380 8412 17382
rect 8468 17380 8492 17382
rect 8548 17380 8572 17382
rect 8628 17380 8652 17382
rect 8708 17380 8714 17382
rect 8406 17371 8714 17380
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 7746 16892 8054 16901
rect 7746 16890 7752 16892
rect 7808 16890 7832 16892
rect 7888 16890 7912 16892
rect 7968 16890 7992 16892
rect 8048 16890 8054 16892
rect 7808 16838 7810 16890
rect 7990 16838 7992 16890
rect 7746 16836 7752 16838
rect 7808 16836 7832 16838
rect 7888 16836 7912 16838
rect 7968 16836 7992 16838
rect 8048 16836 8054 16838
rect 7746 16827 8054 16836
rect 8128 16726 8156 16934
rect 8116 16720 8168 16726
rect 8312 16674 8340 17138
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16794 8524 17070
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8116 16662 8168 16668
rect 7300 16510 7420 16538
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14618 6500 14758
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6932 14498 6960 14962
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14618 7052 14758
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6748 14414 6776 14486
rect 6932 14470 7052 14498
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 14006 6592 14214
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 5632 13320 5684 13326
rect 4908 13246 5028 13274
rect 5632 13262 5684 13268
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12986 4936 13126
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4540 12702 4844 12730
rect 4540 11762 4568 12702
rect 5000 12458 5028 13246
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5276 12481 5304 13194
rect 4724 12430 5028 12458
rect 5262 12472 5318 12481
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 10810 4476 11086
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4540 9994 4568 11698
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4724 9586 4752 12430
rect 5644 12442 5672 13262
rect 6196 12986 6224 13330
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5262 12407 5318 12416
rect 5632 12436 5684 12442
rect 5276 12345 5304 12407
rect 5632 12378 5684 12384
rect 6000 12368 6052 12374
rect 5262 12336 5318 12345
rect 6000 12310 6052 12316
rect 5262 12271 5318 12280
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5000 10674 5028 11766
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5000 10266 5028 10610
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4724 8838 4752 9522
rect 4816 9382 4844 9862
rect 5092 9518 5120 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 9994 5212 10406
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 6012 9654 6040 12310
rect 6196 11762 6224 12922
rect 6288 12374 6316 13806
rect 6380 13530 6408 13806
rect 7024 13734 7052 14470
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6380 12714 6408 13466
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6288 11898 6316 12038
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6380 11762 6408 12650
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6472 10674 6500 12174
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11830 6960 12038
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 11354 6684 11630
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6656 10130 6684 11154
rect 7024 11150 7052 13670
rect 7116 13530 7144 14418
rect 7208 14346 7236 15098
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7300 11218 7328 16510
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7392 16046 7420 16390
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7484 15706 7512 16118
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7668 14550 7696 16390
rect 7746 15804 8054 15813
rect 7746 15802 7752 15804
rect 7808 15802 7832 15804
rect 7888 15802 7912 15804
rect 7968 15802 7992 15804
rect 8048 15802 8054 15804
rect 7808 15750 7810 15802
rect 7990 15750 7992 15802
rect 7746 15748 7752 15750
rect 7808 15748 7832 15750
rect 7888 15748 7912 15750
rect 7968 15748 7992 15750
rect 8048 15748 8054 15750
rect 7746 15739 8054 15748
rect 8128 15638 8156 16662
rect 8220 16646 8340 16674
rect 8220 16250 8248 16646
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8312 16250 8340 16526
rect 8406 16348 8714 16357
rect 8406 16346 8412 16348
rect 8468 16346 8492 16348
rect 8548 16346 8572 16348
rect 8628 16346 8652 16348
rect 8708 16346 8714 16348
rect 8468 16294 8470 16346
rect 8650 16294 8652 16346
rect 8406 16292 8412 16294
rect 8468 16292 8492 16294
rect 8548 16292 8572 16294
rect 8628 16292 8652 16294
rect 8708 16292 8714 16294
rect 8406 16283 8714 16292
rect 8772 16250 8800 16730
rect 8956 16658 8984 19654
rect 9036 19440 9088 19446
rect 9036 19382 9088 19388
rect 9048 18222 9076 19382
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8406 15260 8714 15269
rect 8406 15258 8412 15260
rect 8468 15258 8492 15260
rect 8548 15258 8572 15260
rect 8628 15258 8652 15260
rect 8708 15258 8714 15260
rect 8468 15206 8470 15258
rect 8650 15206 8652 15258
rect 8406 15204 8412 15206
rect 8468 15204 8492 15206
rect 8548 15204 8572 15206
rect 8628 15204 8652 15206
rect 8708 15204 8714 15206
rect 8406 15195 8714 15204
rect 7746 14716 8054 14725
rect 7746 14714 7752 14716
rect 7808 14714 7832 14716
rect 7888 14714 7912 14716
rect 7968 14714 7992 14716
rect 8048 14714 8054 14716
rect 7808 14662 7810 14714
rect 7990 14662 7992 14714
rect 7746 14660 7752 14662
rect 7808 14660 7832 14662
rect 7888 14660 7912 14662
rect 7968 14660 7992 14662
rect 8048 14660 8054 14662
rect 7746 14651 8054 14660
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 12986 7512 14350
rect 8406 14172 8714 14181
rect 8406 14170 8412 14172
rect 8468 14170 8492 14172
rect 8548 14170 8572 14172
rect 8628 14170 8652 14172
rect 8708 14170 8714 14172
rect 8468 14118 8470 14170
rect 8650 14118 8652 14170
rect 8406 14116 8412 14118
rect 8468 14116 8492 14118
rect 8548 14116 8572 14118
rect 8628 14116 8652 14118
rect 8708 14116 8714 14118
rect 8406 14107 8714 14116
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 7746 13628 8054 13637
rect 7746 13626 7752 13628
rect 7808 13626 7832 13628
rect 7888 13626 7912 13628
rect 7968 13626 7992 13628
rect 8048 13626 8054 13628
rect 7808 13574 7810 13626
rect 7990 13574 7992 13626
rect 7746 13572 7752 13574
rect 7808 13572 7832 13574
rect 7888 13572 7912 13574
rect 7968 13572 7992 13574
rect 8048 13572 8054 13574
rect 7746 13563 8054 13572
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7668 12850 7696 13398
rect 8128 13394 8156 13670
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12986 8156 13126
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8312 12918 8340 13874
rect 8772 13734 8800 15574
rect 8956 15502 8984 16594
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 9048 13326 9076 14214
rect 9140 14006 9168 14214
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9036 13320 9088 13326
rect 9232 13274 9260 19926
rect 9324 19854 9352 21714
rect 9876 19854 9904 21714
rect 10428 19854 10456 21714
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 10416 19848 10468 19854
rect 10980 19836 11008 21714
rect 11532 19854 11560 21714
rect 12084 19854 12112 21714
rect 12277 20156 12585 20165
rect 12277 20154 12283 20156
rect 12339 20154 12363 20156
rect 12419 20154 12443 20156
rect 12499 20154 12523 20156
rect 12579 20154 12585 20156
rect 12339 20102 12341 20154
rect 12521 20102 12523 20154
rect 12277 20100 12283 20102
rect 12339 20100 12363 20102
rect 12419 20100 12443 20102
rect 12499 20100 12523 20102
rect 12579 20100 12585 20102
rect 12277 20091 12585 20100
rect 12636 19854 12664 21714
rect 13188 19922 13216 21714
rect 13740 20074 13768 21714
rect 13740 20058 13860 20074
rect 13740 20052 13872 20058
rect 13740 20046 13820 20052
rect 13820 19994 13872 20000
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 14292 19854 14320 21714
rect 11060 19848 11112 19854
rect 10980 19808 11060 19836
rect 10416 19790 10468 19796
rect 11060 19790 11112 19796
rect 11520 19848 11572 19854
rect 12072 19848 12124 19854
rect 11520 19790 11572 19796
rect 11716 19774 11928 19802
rect 12072 19790 12124 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14556 19848 14608 19854
rect 15120 19836 15148 21814
rect 15382 21714 15438 22514
rect 15934 21714 15990 22514
rect 16486 21714 16542 22514
rect 17038 21714 17094 22514
rect 17590 21714 17646 22514
rect 18142 21714 18198 22514
rect 18694 21714 18750 22514
rect 15396 19854 15424 21714
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15200 19848 15252 19854
rect 15120 19808 15200 19836
rect 14556 19790 14608 19796
rect 15200 19790 15252 19796
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9324 18358 9352 18906
rect 9416 18698 9444 19654
rect 10152 19514 10180 19654
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9416 18426 9444 18634
rect 9692 18426 9720 19246
rect 9784 18834 9812 19314
rect 10152 18970 10180 19314
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18970 10272 19110
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9876 18426 9904 18702
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 16250 9536 16526
rect 9692 16250 9720 18090
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9876 15706 9904 16118
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9968 15638 9996 18226
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17882 10088 18022
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10152 17678 10180 18770
rect 10336 18290 10364 19450
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10428 18222 10456 18566
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 16794 10180 17614
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 10428 15094 10456 18158
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10704 16114 10732 16730
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10416 15088 10468 15094
rect 10416 15030 10468 15036
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 14618 9904 14894
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10520 14618 10548 14758
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 9036 13262 9088 13268
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8406 13084 8714 13093
rect 8406 13082 8412 13084
rect 8468 13082 8492 13084
rect 8548 13082 8572 13084
rect 8628 13082 8652 13084
rect 8708 13082 8714 13084
rect 8468 13030 8470 13082
rect 8650 13030 8652 13082
rect 8406 13028 8412 13030
rect 8468 13028 8492 13030
rect 8548 13028 8572 13030
rect 8628 13028 8652 13030
rect 8708 13028 8714 13030
rect 8406 13019 8714 13028
rect 8956 12918 8984 13126
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12442 7696 12786
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 7746 12540 8054 12549
rect 7746 12538 7752 12540
rect 7808 12538 7832 12540
rect 7888 12538 7912 12540
rect 7968 12538 7992 12540
rect 8048 12538 8054 12540
rect 7808 12486 7810 12538
rect 7990 12486 7992 12538
rect 7746 12484 7752 12486
rect 7808 12484 7832 12486
rect 7888 12484 7912 12486
rect 7968 12484 7992 12486
rect 8048 12484 8054 12486
rect 7746 12475 8054 12484
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11898 8156 12174
rect 8406 11996 8714 12005
rect 8406 11994 8412 11996
rect 8468 11994 8492 11996
rect 8548 11994 8572 11996
rect 8628 11994 8652 11996
rect 8708 11994 8714 11996
rect 8468 11942 8470 11994
rect 8650 11942 8652 11994
rect 8406 11940 8412 11942
rect 8468 11940 8492 11942
rect 8548 11940 8572 11942
rect 8628 11940 8652 11942
rect 8708 11940 8714 11942
rect 8406 11931 8714 11940
rect 8956 11898 8984 12718
rect 9048 12374 9076 13262
rect 9140 13246 9260 13274
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 7746 11452 8054 11461
rect 7746 11450 7752 11452
rect 7808 11450 7832 11452
rect 7888 11450 7912 11452
rect 7968 11450 7992 11452
rect 8048 11450 8054 11452
rect 7808 11398 7810 11450
rect 7990 11398 7992 11450
rect 7746 11396 7752 11398
rect 7808 11396 7832 11398
rect 7888 11396 7912 11398
rect 7968 11396 7992 11398
rect 8048 11396 8054 11398
rect 7746 11387 8054 11396
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 5000 7886 5028 8910
rect 5092 8616 5120 9318
rect 6012 8634 6040 9590
rect 6472 8906 6500 9862
rect 6656 9518 6684 10066
rect 6840 9586 6868 10610
rect 7300 10130 7328 11154
rect 8406 10908 8714 10917
rect 8406 10906 8412 10908
rect 8468 10906 8492 10908
rect 8548 10906 8572 10908
rect 8628 10906 8652 10908
rect 8708 10906 8714 10908
rect 8468 10854 8470 10906
rect 8650 10854 8652 10906
rect 8406 10852 8412 10854
rect 8468 10852 8492 10854
rect 8548 10852 8572 10854
rect 8628 10852 8652 10854
rect 8708 10852 8714 10854
rect 8406 10843 8714 10852
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7484 9926 7512 10610
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 10266 7604 10406
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 7024 9518 7052 9862
rect 7668 9586 7696 10542
rect 7746 10364 8054 10373
rect 7746 10362 7752 10364
rect 7808 10362 7832 10364
rect 7888 10362 7912 10364
rect 7968 10362 7992 10364
rect 8048 10362 8054 10364
rect 7808 10310 7810 10362
rect 7990 10310 7992 10362
rect 7746 10308 7752 10310
rect 7808 10308 7832 10310
rect 7888 10308 7912 10310
rect 7968 10308 7992 10310
rect 8048 10308 8054 10310
rect 7746 10299 8054 10308
rect 9048 10062 9076 12310
rect 9140 11898 9168 13246
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12832 9260 13126
rect 9232 12804 9444 12832
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9324 11762 9352 11834
rect 9416 11762 9444 12804
rect 9772 12640 9824 12646
rect 9692 12588 9772 12594
rect 9692 12582 9824 12588
rect 9692 12566 9812 12582
rect 9692 11762 9720 12566
rect 9770 12336 9826 12345
rect 9770 12271 9772 12280
rect 9824 12271 9826 12280
rect 9772 12242 9824 12248
rect 9876 11898 9904 14554
rect 10704 14482 10732 16050
rect 10796 15570 10824 19654
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11072 18850 11100 19382
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10980 18834 11100 18850
rect 10968 18828 11100 18834
rect 11020 18822 11100 18828
rect 10968 18770 11020 18776
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11072 17066 11100 18158
rect 11164 18154 11192 19246
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17338 11192 17546
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11256 16130 11284 19654
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11348 18086 11376 19314
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11624 18766 11652 19110
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 17270 11376 18022
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11716 16130 11744 19774
rect 11900 19718 11928 19774
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 11256 16102 11468 16130
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 15026 10824 15506
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10888 14822 10916 15982
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15706 11192 15846
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14618 10916 14758
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13326 10088 13670
rect 10704 13394 10732 14418
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10888 14074 10916 14282
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10980 13938 11008 15574
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10980 13818 11008 13874
rect 10980 13790 11192 13818
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10060 12782 10088 13262
rect 10244 12986 10272 13262
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11072 12986 11100 13194
rect 11164 13002 11192 13790
rect 11164 12986 11376 13002
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11152 12980 11376 12986
rect 11204 12974 11376 12980
rect 11152 12922 11204 12928
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9312 11756 9364 11762
rect 9232 11716 9312 11744
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7668 9178 7696 9522
rect 8312 9450 8340 9998
rect 9232 9994 9260 11716
rect 9312 11698 9364 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8406 9820 8714 9829
rect 8406 9818 8412 9820
rect 8468 9818 8492 9820
rect 8548 9818 8572 9820
rect 8628 9818 8652 9820
rect 8708 9818 8714 9820
rect 8468 9766 8470 9818
rect 8650 9766 8652 9818
rect 8406 9764 8412 9766
rect 8468 9764 8492 9766
rect 8548 9764 8572 9766
rect 8628 9764 8652 9766
rect 8708 9764 8714 9766
rect 8406 9755 8714 9764
rect 8956 9654 8984 9862
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 7746 9276 8054 9285
rect 7746 9274 7752 9276
rect 7808 9274 7832 9276
rect 7888 9274 7912 9276
rect 7968 9274 7992 9276
rect 8048 9274 8054 9276
rect 7808 9222 7810 9274
rect 7990 9222 7992 9274
rect 7746 9220 7752 9222
rect 7808 9220 7832 9222
rect 7888 9220 7912 9222
rect 7968 9220 7992 9222
rect 8048 9220 8054 9222
rect 7746 9211 8054 9220
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 5172 8628 5224 8634
rect 5092 8588 5172 8616
rect 5092 8294 5120 8588
rect 5172 8570 5224 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7970 5120 8230
rect 5552 8090 5580 8502
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5092 7942 5212 7970
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 7154 3188 7346
rect 3068 7126 3188 7154
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2608 5778 2636 6802
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2700 5574 2728 6666
rect 3068 6458 3096 7126
rect 3215 7100 3523 7109
rect 3215 7098 3221 7100
rect 3277 7098 3301 7100
rect 3357 7098 3381 7100
rect 3437 7098 3461 7100
rect 3517 7098 3523 7100
rect 3277 7046 3279 7098
rect 3459 7046 3461 7098
rect 3215 7044 3221 7046
rect 3277 7044 3301 7046
rect 3357 7044 3381 7046
rect 3437 7044 3461 7046
rect 3517 7044 3523 7046
rect 3215 7035 3523 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6458 3188 6598
rect 3875 6556 4183 6565
rect 3875 6554 3881 6556
rect 3937 6554 3961 6556
rect 4017 6554 4041 6556
rect 4097 6554 4121 6556
rect 4177 6554 4183 6556
rect 3937 6502 3939 6554
rect 4119 6502 4121 6554
rect 3875 6500 3881 6502
rect 3937 6500 3961 6502
rect 4017 6500 4041 6502
rect 4097 6500 4121 6502
rect 4177 6500 4183 6502
rect 3875 6491 4183 6500
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3215 6012 3523 6021
rect 3215 6010 3221 6012
rect 3277 6010 3301 6012
rect 3357 6010 3381 6012
rect 3437 6010 3461 6012
rect 3517 6010 3523 6012
rect 3277 5958 3279 6010
rect 3459 5958 3461 6010
rect 3215 5956 3221 5958
rect 3277 5956 3301 5958
rect 3357 5956 3381 5958
rect 3437 5956 3461 5958
rect 3517 5956 3523 5958
rect 3215 5947 3523 5956
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 1768 5092 1820 5098
rect 1768 5034 1820 5040
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 1780 4690 1808 5034
rect 2516 4690 2544 5510
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2700 4146 2728 5510
rect 2976 5370 3004 5646
rect 3804 5642 3832 6190
rect 4264 5778 4292 6938
rect 4356 6662 4384 7822
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7546 4660 7686
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 5000 7002 5028 7822
rect 5092 7546 5120 7822
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4632 5710 4660 6054
rect 4620 5704 4672 5710
rect 5000 5692 5028 6938
rect 5184 6866 5212 7942
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5184 6458 5212 6802
rect 5552 6798 5580 7346
rect 6012 7342 6040 8230
rect 6656 7818 6684 8978
rect 9232 8974 9260 9318
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7024 8634 7052 8842
rect 8406 8732 8714 8741
rect 8406 8730 8412 8732
rect 8468 8730 8492 8732
rect 8548 8730 8572 8732
rect 8628 8730 8652 8732
rect 8708 8730 8714 8732
rect 8468 8678 8470 8730
rect 8650 8678 8652 8730
rect 8406 8676 8412 8678
rect 8468 8676 8492 8678
rect 8548 8676 8572 8678
rect 8628 8676 8652 8678
rect 8708 8676 8714 8678
rect 8406 8667 8714 8676
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 8242 8340 8434
rect 8220 8214 8340 8242
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 7746 8188 8054 8197
rect 7746 8186 7752 8188
rect 7808 8186 7832 8188
rect 7888 8186 7912 8188
rect 7968 8186 7992 8188
rect 8048 8186 8054 8188
rect 7808 8134 7810 8186
rect 7990 8134 7992 8186
rect 7746 8132 7752 8134
rect 7808 8132 7832 8134
rect 7888 8132 7912 8134
rect 7968 8132 7992 8134
rect 8048 8132 8054 8134
rect 7746 8123 8054 8132
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5710 5304 6190
rect 5172 5704 5224 5710
rect 5000 5664 5172 5692
rect 4620 5646 4672 5652
rect 5172 5646 5224 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3215 4924 3523 4933
rect 3215 4922 3221 4924
rect 3277 4922 3301 4924
rect 3357 4922 3381 4924
rect 3437 4922 3461 4924
rect 3517 4922 3523 4924
rect 3277 4870 3279 4922
rect 3459 4870 3461 4922
rect 3215 4868 3221 4870
rect 3277 4868 3301 4870
rect 3357 4868 3381 4870
rect 3437 4868 3461 4870
rect 3517 4868 3523 4870
rect 3215 4859 3523 4868
rect 3804 4826 3832 5578
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 3875 5468 4183 5477
rect 3875 5466 3881 5468
rect 3937 5466 3961 5468
rect 4017 5466 4041 5468
rect 4097 5466 4121 5468
rect 4177 5466 4183 5468
rect 3937 5414 3939 5466
rect 4119 5414 4121 5466
rect 3875 5412 3881 5414
rect 3937 5412 3961 5414
rect 4017 5412 4041 5414
rect 4097 5412 4121 5414
rect 4177 5412 4183 5414
rect 3875 5403 4183 5412
rect 4908 5370 4936 5510
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 5368 5166 5396 5578
rect 5460 5166 5488 6598
rect 7024 6322 7052 7754
rect 7116 7546 7144 7822
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7668 6390 7696 7958
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7546 7788 7686
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7944 7274 7972 7890
rect 8220 7750 8248 8214
rect 8772 7954 8800 8230
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7546 8248 7686
rect 8406 7644 8714 7653
rect 8406 7642 8412 7644
rect 8468 7642 8492 7644
rect 8548 7642 8572 7644
rect 8628 7642 8652 7644
rect 8708 7642 8714 7644
rect 8468 7590 8470 7642
rect 8650 7590 8652 7642
rect 8406 7588 8412 7590
rect 8468 7588 8492 7590
rect 8548 7588 8572 7590
rect 8628 7588 8652 7590
rect 8708 7588 8714 7590
rect 8406 7579 8714 7588
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7746 7100 8054 7109
rect 7746 7098 7752 7100
rect 7808 7098 7832 7100
rect 7888 7098 7912 7100
rect 7968 7098 7992 7100
rect 8048 7098 8054 7100
rect 7808 7046 7810 7098
rect 7990 7046 7992 7098
rect 7746 7044 7752 7046
rect 7808 7044 7832 7046
rect 7888 7044 7912 7046
rect 7968 7044 7992 7046
rect 8048 7044 8054 7046
rect 7746 7035 8054 7044
rect 8956 7002 8984 7414
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8406 6556 8714 6565
rect 8406 6554 8412 6556
rect 8468 6554 8492 6556
rect 8548 6554 8572 6556
rect 8628 6554 8652 6556
rect 8708 6554 8714 6556
rect 8468 6502 8470 6554
rect 8650 6502 8652 6554
rect 8406 6500 8412 6502
rect 8468 6500 8492 6502
rect 8548 6500 8572 6502
rect 8628 6500 8652 6502
rect 8708 6500 8714 6502
rect 8406 6491 8714 6500
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6932 5370 6960 5578
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 4172 4826 4200 5102
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4264 4690 4292 5102
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 5460 4622 5488 5102
rect 5736 4826 5764 5238
rect 7024 5234 7052 6258
rect 7746 6012 8054 6021
rect 7746 6010 7752 6012
rect 7808 6010 7832 6012
rect 7888 6010 7912 6012
rect 7968 6010 7992 6012
rect 8048 6010 8054 6012
rect 7808 5958 7810 6010
rect 7990 5958 7992 6010
rect 7746 5956 7752 5958
rect 7808 5956 7832 5958
rect 7888 5956 7912 5958
rect 7968 5956 7992 5958
rect 8048 5956 8054 5958
rect 7746 5947 8054 5956
rect 8772 5846 8800 6598
rect 9232 6236 9260 8910
rect 9324 8566 9352 10542
rect 9416 9654 9444 11562
rect 9784 11354 9812 11698
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 11218 9904 11834
rect 10612 11218 10640 12718
rect 11256 12442 11284 12786
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10810 10456 10950
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10612 10266 10640 11154
rect 10796 11150 10824 11494
rect 11072 11257 11100 12106
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11286 11192 12038
rect 11152 11280 11204 11286
rect 11058 11248 11114 11257
rect 11152 11222 11204 11228
rect 11058 11183 11114 11192
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10810 11100 11018
rect 11164 10810 11192 11086
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 10968 8968 11020 8974
rect 11072 8956 11100 10610
rect 11256 10606 11284 10950
rect 11348 10674 11376 12974
rect 11440 12170 11468 16102
rect 11624 16102 11744 16130
rect 11808 16130 11836 19654
rect 12937 19612 13245 19621
rect 12937 19610 12943 19612
rect 12999 19610 13023 19612
rect 13079 19610 13103 19612
rect 13159 19610 13183 19612
rect 13239 19610 13245 19612
rect 12999 19558 13001 19610
rect 13181 19558 13183 19610
rect 12937 19556 12943 19558
rect 12999 19556 13023 19558
rect 13079 19556 13103 19558
rect 13159 19556 13183 19558
rect 13239 19556 13245 19558
rect 12937 19547 13245 19556
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12277 19068 12585 19077
rect 12277 19066 12283 19068
rect 12339 19066 12363 19068
rect 12419 19066 12443 19068
rect 12499 19066 12523 19068
rect 12579 19066 12585 19068
rect 12339 19014 12341 19066
rect 12521 19014 12523 19066
rect 12277 19012 12283 19014
rect 12339 19012 12363 19014
rect 12419 19012 12443 19014
rect 12499 19012 12523 19014
rect 12579 19012 12585 19014
rect 12277 19003 12585 19012
rect 12636 18970 12664 19246
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18358 12112 18566
rect 12937 18524 13245 18533
rect 12937 18522 12943 18524
rect 12999 18522 13023 18524
rect 13079 18522 13103 18524
rect 13159 18522 13183 18524
rect 13239 18522 13245 18524
rect 12999 18470 13001 18522
rect 13181 18470 13183 18522
rect 12937 18468 12943 18470
rect 12999 18468 13023 18470
rect 13079 18468 13103 18470
rect 13159 18468 13183 18470
rect 13239 18468 13245 18470
rect 12937 18459 13245 18468
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11992 17134 12020 18158
rect 12277 17980 12585 17989
rect 12277 17978 12283 17980
rect 12339 17978 12363 17980
rect 12419 17978 12443 17980
rect 12499 17978 12523 17980
rect 12579 17978 12585 17980
rect 12339 17926 12341 17978
rect 12521 17926 12523 17978
rect 12277 17924 12283 17926
rect 12339 17924 12363 17926
rect 12419 17924 12443 17926
rect 12499 17924 12523 17926
rect 12579 17924 12585 17926
rect 12277 17915 12585 17924
rect 13280 17746 13308 18770
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 12360 17338 12388 17682
rect 13372 17678 13400 18022
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12820 17338 12848 17478
rect 12937 17436 13245 17445
rect 12937 17434 12943 17436
rect 12999 17434 13023 17436
rect 13079 17434 13103 17436
rect 13159 17434 13183 17436
rect 13239 17434 13245 17436
rect 12999 17382 13001 17434
rect 13181 17382 13183 17434
rect 12937 17380 12943 17382
rect 12999 17380 13023 17382
rect 13079 17380 13103 17382
rect 13159 17380 13183 17382
rect 13239 17380 13245 17382
rect 12937 17371 13245 17380
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 12277 16892 12585 16901
rect 12277 16890 12283 16892
rect 12339 16890 12363 16892
rect 12419 16890 12443 16892
rect 12499 16890 12523 16892
rect 12579 16890 12585 16892
rect 12339 16838 12341 16890
rect 12521 16838 12523 16890
rect 12277 16836 12283 16838
rect 12339 16836 12363 16838
rect 12419 16836 12443 16838
rect 12499 16836 12523 16838
rect 12579 16836 12585 16838
rect 12277 16827 12585 16836
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12072 16176 12124 16182
rect 11808 16102 11928 16130
rect 12072 16118 12124 16124
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11532 12238 11560 15302
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11532 11914 11560 12174
rect 11440 11898 11560 11914
rect 11440 11892 11572 11898
rect 11440 11886 11520 11892
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9722 11192 10066
rect 11256 10062 11284 10542
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11440 9874 11468 11886
rect 11520 11834 11572 11840
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11256 9846 11468 9874
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11256 9586 11284 9846
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11532 9518 11560 11630
rect 11624 11218 11652 16102
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14074 11744 14894
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 14074 11836 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12986 11836 13194
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11716 10266 11744 10610
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11164 9178 11192 9386
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9178 11284 9318
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11020 8928 11100 8956
rect 10968 8910 11020 8916
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9416 7886 9444 8910
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9876 8090 9904 8502
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 10152 7750 10180 8774
rect 10704 8634 10732 8774
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11072 7886 11100 8928
rect 11532 8430 11560 9454
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11532 8090 11560 8366
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 9692 7546 9720 7686
rect 10152 7546 10180 7686
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10336 7478 10364 7822
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7546 10456 7686
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 11532 7410 11560 8026
rect 11624 7886 11652 9930
rect 11716 9518 11744 9998
rect 11900 9654 11928 16102
rect 12084 15706 12112 16118
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12176 13512 12204 16458
rect 12820 16250 12848 17138
rect 12937 16348 13245 16357
rect 12937 16346 12943 16348
rect 12999 16346 13023 16348
rect 13079 16346 13103 16348
rect 13159 16346 13183 16348
rect 13239 16346 13245 16348
rect 12999 16294 13001 16346
rect 13181 16294 13183 16346
rect 12937 16292 12943 16294
rect 12999 16292 13023 16294
rect 13079 16292 13103 16294
rect 13159 16292 13183 16294
rect 13239 16292 13245 16294
rect 12937 16283 13245 16292
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12277 15804 12585 15813
rect 12277 15802 12283 15804
rect 12339 15802 12363 15804
rect 12419 15802 12443 15804
rect 12499 15802 12523 15804
rect 12579 15802 12585 15804
rect 12339 15750 12341 15802
rect 12521 15750 12523 15802
rect 12277 15748 12283 15750
rect 12339 15748 12363 15750
rect 12419 15748 12443 15750
rect 12499 15748 12523 15750
rect 12579 15748 12585 15750
rect 12277 15739 12585 15748
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12452 15162 12480 15370
rect 12937 15260 13245 15269
rect 12937 15258 12943 15260
rect 12999 15258 13023 15260
rect 13079 15258 13103 15260
rect 13159 15258 13183 15260
rect 13239 15258 13245 15260
rect 12999 15206 13001 15258
rect 13181 15206 13183 15258
rect 12937 15204 12943 15206
rect 12999 15204 13023 15206
rect 13079 15204 13103 15206
rect 13159 15204 13183 15206
rect 13239 15204 13245 15206
rect 12937 15195 13245 15204
rect 13464 15162 13492 19654
rect 13648 19446 13676 19654
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13740 18834 13768 19654
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 16998 13584 18566
rect 13648 17202 13676 18634
rect 13740 18426 13768 18770
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 17338 13768 17478
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13556 15042 13584 16934
rect 13648 15570 13676 17138
rect 14016 17134 14044 19654
rect 14200 18834 14228 19654
rect 14384 19514 14412 19790
rect 14568 19514 14596 19790
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14568 18766 14596 19450
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 15120 17678 15148 19654
rect 15396 19378 15424 19654
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15212 18426 15240 18634
rect 15304 18426 15332 19110
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15396 18154 15424 19110
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14936 16046 14964 17002
rect 15120 16658 15148 17614
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15706 13860 15846
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 13464 15014 13584 15042
rect 13464 14958 13492 15014
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12277 14716 12585 14725
rect 12277 14714 12283 14716
rect 12339 14714 12363 14716
rect 12419 14714 12443 14716
rect 12499 14714 12523 14716
rect 12579 14714 12585 14716
rect 12339 14662 12341 14714
rect 12521 14662 12523 14714
rect 12277 14660 12283 14662
rect 12339 14660 12363 14662
rect 12419 14660 12443 14662
rect 12499 14660 12523 14662
rect 12579 14660 12585 14662
rect 12277 14651 12585 14660
rect 13556 14618 13584 14758
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13648 14482 13676 15506
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 13924 15026 13952 15302
rect 14292 15026 14320 15302
rect 14476 15026 14504 15506
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14618 13860 14758
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 12820 13870 12848 14418
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 12937 14172 13245 14181
rect 12937 14170 12943 14172
rect 12999 14170 13023 14172
rect 13079 14170 13103 14172
rect 13159 14170 13183 14172
rect 13239 14170 13245 14172
rect 12999 14118 13001 14170
rect 13181 14118 13183 14170
rect 12937 14116 12943 14118
rect 12999 14116 13023 14118
rect 13079 14116 13103 14118
rect 13159 14116 13183 14118
rect 13239 14116 13245 14118
rect 12937 14107 13245 14116
rect 13280 13870 13308 14214
rect 13648 14090 13676 14418
rect 13556 14074 13676 14090
rect 13544 14068 13676 14074
rect 13596 14062 13676 14068
rect 13544 14010 13596 14016
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 12277 13628 12585 13637
rect 12277 13626 12283 13628
rect 12339 13626 12363 13628
rect 12419 13626 12443 13628
rect 12499 13626 12523 13628
rect 12579 13626 12585 13628
rect 12339 13574 12341 13626
rect 12521 13574 12523 13626
rect 12277 13572 12283 13574
rect 12339 13572 12363 13574
rect 12419 13572 12443 13574
rect 12499 13572 12523 13574
rect 12579 13572 12585 13574
rect 12277 13563 12585 13572
rect 12820 13530 12848 13806
rect 12808 13524 12860 13530
rect 12176 13484 12296 13512
rect 12268 13410 12296 13484
rect 12808 13466 12860 13472
rect 12268 13382 12664 13410
rect 12636 12918 12664 13382
rect 12937 13084 13245 13093
rect 12937 13082 12943 13084
rect 12999 13082 13023 13084
rect 13079 13082 13103 13084
rect 13159 13082 13183 13084
rect 13239 13082 13245 13084
rect 12999 13030 13001 13082
rect 13181 13030 13183 13082
rect 12937 13028 12943 13030
rect 12999 13028 13023 13030
rect 13079 13028 13103 13030
rect 13159 13028 13183 13030
rect 13239 13028 13245 13030
rect 12937 13019 13245 13028
rect 14384 12986 14412 14418
rect 14936 13938 14964 15982
rect 15396 15502 15424 16934
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15396 14958 15424 15438
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15304 14074 15332 14282
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12277 12540 12585 12549
rect 12277 12538 12283 12540
rect 12339 12538 12363 12540
rect 12419 12538 12443 12540
rect 12499 12538 12523 12540
rect 12579 12538 12585 12540
rect 12339 12486 12341 12538
rect 12521 12486 12523 12538
rect 12277 12484 12283 12486
rect 12339 12484 12363 12486
rect 12419 12484 12443 12486
rect 12499 12484 12523 12486
rect 12579 12484 12585 12486
rect 12277 12475 12585 12484
rect 12636 12434 12664 12854
rect 12636 12406 12848 12434
rect 12820 12345 12848 12406
rect 12806 12336 12862 12345
rect 12806 12271 12862 12280
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12176 11354 12204 11766
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12277 11452 12585 11461
rect 12277 11450 12283 11452
rect 12339 11450 12363 11452
rect 12419 11450 12443 11452
rect 12499 11450 12523 11452
rect 12579 11450 12585 11452
rect 12339 11398 12341 11450
rect 12521 11398 12523 11450
rect 12277 11396 12283 11398
rect 12339 11396 12363 11398
rect 12419 11396 12443 11398
rect 12499 11396 12523 11398
rect 12579 11396 12585 11398
rect 12277 11387 12585 11396
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12636 11218 12664 11494
rect 12728 11286 12756 12038
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12452 10606 12480 11154
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12277 10364 12585 10373
rect 12277 10362 12283 10364
rect 12339 10362 12363 10364
rect 12419 10362 12443 10364
rect 12499 10362 12523 10364
rect 12579 10362 12585 10364
rect 12339 10310 12341 10362
rect 12521 10310 12523 10362
rect 12277 10308 12283 10310
rect 12339 10308 12363 10310
rect 12419 10308 12443 10310
rect 12499 10308 12523 10310
rect 12579 10308 12585 10310
rect 12277 10299 12585 10308
rect 12636 10266 12664 11154
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10674 12756 10950
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 12636 9586 12664 10202
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 11716 8634 11744 9454
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 8634 12020 9318
rect 12277 9276 12585 9285
rect 12277 9274 12283 9276
rect 12339 9274 12363 9276
rect 12419 9274 12443 9276
rect 12499 9274 12523 9276
rect 12579 9274 12585 9276
rect 12339 9222 12341 9274
rect 12521 9222 12523 9274
rect 12277 9220 12283 9222
rect 12339 9220 12363 9222
rect 12419 9220 12443 9222
rect 12499 9220 12523 9222
rect 12579 9220 12585 9222
rect 12277 9211 12585 9220
rect 12728 9178 12756 9454
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12820 8430 12848 12271
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 12937 11996 13245 12005
rect 12937 11994 12943 11996
rect 12999 11994 13023 11996
rect 13079 11994 13103 11996
rect 13159 11994 13183 11996
rect 13239 11994 13245 11996
rect 12999 11942 13001 11994
rect 13181 11942 13183 11994
rect 12937 11940 12943 11942
rect 12999 11940 13023 11942
rect 13079 11940 13103 11942
rect 13159 11940 13183 11942
rect 13239 11940 13245 11942
rect 12937 11931 13245 11940
rect 13832 11898 13860 12174
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11354 12940 11494
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 13096 11150 13124 11834
rect 14200 11762 14228 12038
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 13372 11354 13400 11698
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12937 10908 13245 10917
rect 12937 10906 12943 10908
rect 12999 10906 13023 10908
rect 13079 10906 13103 10908
rect 13159 10906 13183 10908
rect 13239 10906 13245 10908
rect 12999 10854 13001 10906
rect 13181 10854 13183 10906
rect 12937 10852 12943 10854
rect 12999 10852 13023 10854
rect 13079 10852 13103 10854
rect 13159 10852 13183 10854
rect 13239 10852 13245 10854
rect 12937 10843 13245 10852
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 12937 9820 13245 9829
rect 12937 9818 12943 9820
rect 12999 9818 13023 9820
rect 13079 9818 13103 9820
rect 13159 9818 13183 9820
rect 13239 9818 13245 9820
rect 12999 9766 13001 9818
rect 13181 9766 13183 9818
rect 12937 9764 12943 9766
rect 12999 9764 13023 9766
rect 13079 9764 13103 9766
rect 13159 9764 13183 9766
rect 13239 9764 13245 9766
rect 12937 9755 13245 9764
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9178 13400 9386
rect 13648 9382 13676 9998
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13648 9042 13676 9318
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13832 8974 13860 9862
rect 13924 9518 13952 10474
rect 14292 10130 14320 12174
rect 14660 12170 14688 13806
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14660 11694 14688 12106
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14936 11218 14964 13874
rect 15488 12986 15516 19654
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15672 14226 15700 16050
rect 15764 15162 15792 19926
rect 15948 19854 15976 21714
rect 16500 20482 16528 21714
rect 16500 20454 16620 20482
rect 16592 20398 16620 20454
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 17052 20346 17080 21714
rect 17500 20392 17552 20398
rect 17052 20318 17264 20346
rect 17500 20334 17552 20340
rect 16808 20156 17116 20165
rect 16808 20154 16814 20156
rect 16870 20154 16894 20156
rect 16950 20154 16974 20156
rect 17030 20154 17054 20156
rect 17110 20154 17116 20156
rect 16870 20102 16872 20154
rect 17052 20102 17054 20154
rect 16808 20100 16814 20102
rect 16870 20100 16894 20102
rect 16950 20100 16974 20102
rect 17030 20100 17054 20102
rect 17110 20100 17116 20102
rect 16808 20091 17116 20100
rect 17236 19922 17264 20318
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17512 19854 17540 20334
rect 17604 19922 17632 21714
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16580 19848 16632 19854
rect 17500 19848 17552 19854
rect 16580 19790 16632 19796
rect 17130 19816 17186 19825
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 17678 15884 18022
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15856 17338 15884 17478
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16658 15884 16934
rect 16040 16726 16068 17070
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15580 14198 15700 14226
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12306 15332 12582
rect 15580 12434 15608 14198
rect 15764 13938 15792 15098
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15856 13802 15884 16594
rect 16132 15910 16160 17478
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14346 15976 14758
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 16040 14278 16068 14962
rect 16132 14890 16160 15846
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15672 12782 15700 13738
rect 16132 12850 16160 14826
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15488 12406 15608 12434
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15304 11898 15332 12106
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10130 14780 10406
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14292 9654 14320 10066
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14108 9178 14136 9590
rect 14936 9586 14964 11154
rect 15488 10674 15516 12406
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10266 15332 10542
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 12937 8732 13245 8741
rect 12937 8730 12943 8732
rect 12999 8730 13023 8732
rect 13079 8730 13103 8732
rect 13159 8730 13183 8732
rect 13239 8730 13245 8732
rect 12999 8678 13001 8730
rect 13181 8678 13183 8730
rect 12937 8676 12943 8678
rect 12999 8676 13023 8678
rect 13079 8676 13103 8678
rect 13159 8676 13183 8678
rect 13239 8676 13245 8678
rect 12937 8667 13245 8676
rect 13556 8634 13584 8910
rect 14660 8634 14688 9522
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12277 8188 12585 8197
rect 12277 8186 12283 8188
rect 12339 8186 12363 8188
rect 12419 8186 12443 8188
rect 12499 8186 12523 8188
rect 12579 8186 12585 8188
rect 12339 8134 12341 8186
rect 12521 8134 12523 8186
rect 12277 8132 12283 8134
rect 12339 8132 12363 8134
rect 12419 8132 12443 8134
rect 12499 8132 12523 8134
rect 12579 8132 12585 8134
rect 12277 8123 12585 8132
rect 12820 8090 12848 8366
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12912 8022 12940 8434
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 6866 9444 7278
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 10428 6798 10456 7142
rect 10612 7002 10640 7346
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9312 6248 9364 6254
rect 9232 6208 9312 6236
rect 9312 6190 9364 6196
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5914 9260 6054
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8406 5468 8714 5477
rect 8406 5466 8412 5468
rect 8468 5466 8492 5468
rect 8548 5466 8572 5468
rect 8628 5466 8652 5468
rect 8708 5466 8714 5468
rect 8468 5414 8470 5466
rect 8650 5414 8652 5466
rect 8406 5412 8412 5414
rect 8468 5412 8492 5414
rect 8548 5412 8572 5414
rect 8628 5412 8652 5414
rect 8708 5412 8714 5414
rect 8406 5403 8714 5412
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 8772 5166 8800 5782
rect 9232 5710 9260 5850
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9324 5166 9352 6190
rect 9508 5914 9536 6326
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9692 5386 9720 6054
rect 10704 5642 10732 6054
rect 10980 5778 11008 7346
rect 11624 6798 11652 7822
rect 12937 7644 13245 7653
rect 12937 7642 12943 7644
rect 12999 7642 13023 7644
rect 13079 7642 13103 7644
rect 13159 7642 13183 7644
rect 13239 7642 13245 7644
rect 12999 7590 13001 7642
rect 13181 7590 13183 7642
rect 12937 7588 12943 7590
rect 12999 7588 13023 7590
rect 13079 7588 13103 7590
rect 13159 7588 13183 7590
rect 13239 7588 13245 7590
rect 12937 7579 13245 7588
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12277 7100 12585 7109
rect 12277 7098 12283 7100
rect 12339 7098 12363 7100
rect 12419 7098 12443 7100
rect 12499 7098 12523 7100
rect 12579 7098 12585 7100
rect 12339 7046 12341 7098
rect 12521 7046 12523 7098
rect 12277 7044 12283 7046
rect 12339 7044 12363 7046
rect 12419 7044 12443 7046
rect 12499 7044 12523 7046
rect 12579 7044 12585 7046
rect 12277 7035 12585 7044
rect 12912 7002 12940 7414
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13832 6882 13860 8434
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14016 7002 14044 7822
rect 14108 7546 14136 7822
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13740 6866 13860 6882
rect 13728 6860 13860 6866
rect 13780 6854 13860 6860
rect 13728 6802 13780 6808
rect 14108 6798 14136 7278
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 11624 6322 11652 6734
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11808 6254 11836 6598
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5914 11560 6054
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11716 5778 11744 6190
rect 12277 6012 12585 6021
rect 12277 6010 12283 6012
rect 12339 6010 12363 6012
rect 12419 6010 12443 6012
rect 12499 6010 12523 6012
rect 12579 6010 12585 6012
rect 12339 5958 12341 6010
rect 12521 5958 12523 6010
rect 12277 5956 12283 5958
rect 12339 5956 12363 5958
rect 12419 5956 12443 5958
rect 12499 5956 12523 5958
rect 12579 5956 12585 5958
rect 12277 5947 12585 5956
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 9600 5370 9720 5386
rect 9588 5364 9720 5370
rect 9640 5358 9720 5364
rect 9588 5306 9640 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 4826 6224 4966
rect 7746 4924 8054 4933
rect 7746 4922 7752 4924
rect 7808 4922 7832 4924
rect 7888 4922 7912 4924
rect 7968 4922 7992 4924
rect 8048 4922 8054 4924
rect 7808 4870 7810 4922
rect 7990 4870 7992 4922
rect 7746 4868 7752 4870
rect 7808 4868 7832 4870
rect 7888 4868 7912 4870
rect 7968 4868 7992 4870
rect 8048 4868 8054 4870
rect 7746 4859 8054 4868
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 8772 4622 8800 5102
rect 9692 4826 9720 5238
rect 10980 5234 11008 5714
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11624 5370 11652 5646
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11716 5166 11744 5714
rect 11900 5234 11928 5782
rect 12636 5710 12664 6598
rect 12820 6390 12848 6734
rect 12937 6556 13245 6565
rect 12937 6554 12943 6556
rect 12999 6554 13023 6556
rect 13079 6554 13103 6556
rect 13159 6554 13183 6556
rect 13239 6554 13245 6556
rect 12999 6502 13001 6554
rect 13181 6502 13183 6554
rect 12937 6500 12943 6502
rect 12999 6500 13023 6502
rect 13079 6500 13103 6502
rect 13159 6500 13183 6502
rect 13239 6500 13245 6502
rect 12937 6491 13245 6500
rect 12808 6384 12860 6390
rect 12728 6332 12808 6338
rect 12728 6326 12860 6332
rect 12728 6310 12848 6326
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11992 5166 12020 5510
rect 12636 5302 12664 5510
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 12277 4924 12585 4933
rect 12277 4922 12283 4924
rect 12339 4922 12363 4924
rect 12419 4922 12443 4924
rect 12499 4922 12523 4924
rect 12579 4922 12585 4924
rect 12339 4870 12341 4922
rect 12521 4870 12523 4922
rect 12277 4868 12283 4870
rect 12339 4868 12363 4870
rect 12419 4868 12443 4870
rect 12499 4868 12523 4870
rect 12579 4868 12585 4870
rect 12277 4859 12585 4868
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 12728 4622 12756 6310
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5914 12848 6190
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12937 5468 13245 5477
rect 12937 5466 12943 5468
rect 12999 5466 13023 5468
rect 13079 5466 13103 5468
rect 13159 5466 13183 5468
rect 13239 5466 13245 5468
rect 12999 5414 13001 5466
rect 13181 5414 13183 5466
rect 12937 5412 12943 5414
rect 12999 5412 13023 5414
rect 13079 5412 13103 5414
rect 13159 5412 13183 5414
rect 13239 5412 13245 5414
rect 12937 5403 13245 5412
rect 14108 5370 14136 6734
rect 14660 6458 14688 8570
rect 14752 8498 14780 9522
rect 14936 8974 14964 9522
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 7546 14872 7686
rect 14936 7546 14964 7890
rect 15200 7880 15252 7886
rect 15304 7834 15332 8366
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15252 7828 15332 7834
rect 15200 7822 15332 7828
rect 15212 7806 15332 7822
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 15212 7410 15240 7686
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15212 6934 15240 7346
rect 15304 6934 15332 7806
rect 15396 7342 15424 8026
rect 15488 7886 15516 10610
rect 15580 9926 15608 11698
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 8430 15608 9862
rect 15672 9722 15700 12718
rect 15764 11898 15792 12718
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 10198 16068 11698
rect 16224 10810 16252 19654
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16316 18970 16344 19110
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16592 18902 16620 19790
rect 17130 19751 17186 19760
rect 17236 19774 17448 19802
rect 17500 19790 17552 19796
rect 17682 19816 17738 19825
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19514 16712 19654
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16684 18766 16712 19314
rect 16808 19068 17116 19077
rect 16808 19066 16814 19068
rect 16870 19066 16894 19068
rect 16950 19066 16974 19068
rect 17030 19066 17054 19068
rect 17110 19066 17116 19068
rect 16870 19014 16872 19066
rect 17052 19014 17054 19066
rect 16808 19012 16814 19014
rect 16870 19012 16894 19014
rect 16950 19012 16974 19014
rect 17030 19012 17054 19014
rect 17110 19012 17116 19014
rect 16808 19003 17116 19012
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 17202 16620 18566
rect 16684 17746 16712 18702
rect 16776 18222 16804 18770
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16808 17980 17116 17989
rect 16808 17978 16814 17980
rect 16870 17978 16894 17980
rect 16950 17978 16974 17980
rect 17030 17978 17054 17980
rect 17110 17978 17116 17980
rect 16870 17926 16872 17978
rect 17052 17926 17054 17978
rect 16808 17924 16814 17926
rect 16870 17924 16894 17926
rect 16950 17924 16974 17926
rect 17030 17924 17054 17926
rect 17110 17924 17116 17926
rect 16808 17915 17116 17924
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16592 17066 16620 17138
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16592 16250 16620 17002
rect 16684 16658 16712 17682
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 17052 17338 17080 17546
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16808 16892 17116 16901
rect 16808 16890 16814 16892
rect 16870 16890 16894 16892
rect 16950 16890 16974 16892
rect 17030 16890 17054 16892
rect 17110 16890 17116 16892
rect 16870 16838 16872 16890
rect 17052 16838 17054 16890
rect 16808 16836 16814 16838
rect 16870 16836 16894 16838
rect 16950 16836 16974 16838
rect 17030 16836 17054 16838
rect 17110 16836 17116 16838
rect 16808 16827 17116 16836
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 11830 16344 14214
rect 16592 13326 16620 14758
rect 16684 14482 16712 16594
rect 16776 16250 16804 16730
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16808 15804 17116 15813
rect 16808 15802 16814 15804
rect 16870 15802 16894 15804
rect 16950 15802 16974 15804
rect 17030 15802 17054 15804
rect 17110 15802 17116 15804
rect 16870 15750 16872 15802
rect 17052 15750 17054 15802
rect 16808 15748 16814 15750
rect 16870 15748 16894 15750
rect 16950 15748 16974 15750
rect 17030 15748 17054 15750
rect 17110 15748 17116 15750
rect 16808 15739 17116 15748
rect 16808 14716 17116 14725
rect 16808 14714 16814 14716
rect 16870 14714 16894 14716
rect 16950 14714 16974 14716
rect 17030 14714 17054 14716
rect 17110 14714 17116 14716
rect 16870 14662 16872 14714
rect 17052 14662 17054 14714
rect 16808 14660 16814 14662
rect 16870 14660 16894 14662
rect 16950 14660 16974 14662
rect 17030 14660 17054 14662
rect 17110 14660 17116 14662
rect 16808 14651 17116 14660
rect 16948 14612 17000 14618
rect 17144 14600 17172 19751
rect 17236 14770 17264 19774
rect 17420 19718 17448 19774
rect 17682 19751 17738 19760
rect 17696 19718 17724 19751
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17328 16998 17356 19654
rect 17468 19612 17776 19621
rect 17468 19610 17474 19612
rect 17530 19610 17554 19612
rect 17610 19610 17634 19612
rect 17690 19610 17714 19612
rect 17770 19610 17776 19612
rect 17530 19558 17532 19610
rect 17712 19558 17714 19610
rect 17468 19556 17474 19558
rect 17530 19556 17554 19558
rect 17610 19556 17634 19558
rect 17690 19556 17714 19558
rect 17770 19556 17776 19558
rect 17468 19547 17776 19556
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 17420 18970 17448 19382
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17468 18524 17776 18533
rect 17468 18522 17474 18524
rect 17530 18522 17554 18524
rect 17610 18522 17634 18524
rect 17690 18522 17714 18524
rect 17770 18522 17776 18524
rect 17530 18470 17532 18522
rect 17712 18470 17714 18522
rect 17468 18468 17474 18470
rect 17530 18468 17554 18470
rect 17610 18468 17634 18470
rect 17690 18468 17714 18470
rect 17770 18468 17776 18470
rect 17468 18459 17776 18468
rect 17468 17436 17776 17445
rect 17468 17434 17474 17436
rect 17530 17434 17554 17436
rect 17610 17434 17634 17436
rect 17690 17434 17714 17436
rect 17770 17434 17776 17436
rect 17530 17382 17532 17434
rect 17712 17382 17714 17434
rect 17468 17380 17474 17382
rect 17530 17380 17554 17382
rect 17610 17380 17634 17382
rect 17690 17380 17714 17382
rect 17770 17380 17776 17382
rect 17468 17371 17776 17380
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17328 16250 17356 16458
rect 17468 16348 17776 16357
rect 17468 16346 17474 16348
rect 17530 16346 17554 16348
rect 17610 16346 17634 16348
rect 17690 16346 17714 16348
rect 17770 16346 17776 16348
rect 17530 16294 17532 16346
rect 17712 16294 17714 16346
rect 17468 16292 17474 16294
rect 17530 16292 17554 16294
rect 17610 16292 17634 16294
rect 17690 16292 17714 16294
rect 17770 16292 17776 16294
rect 17468 16283 17776 16292
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17468 15260 17776 15269
rect 17468 15258 17474 15260
rect 17530 15258 17554 15260
rect 17610 15258 17634 15260
rect 17690 15258 17714 15260
rect 17770 15258 17776 15260
rect 17530 15206 17532 15258
rect 17712 15206 17714 15258
rect 17468 15204 17474 15206
rect 17530 15204 17554 15206
rect 17610 15204 17634 15206
rect 17690 15204 17714 15206
rect 17770 15204 17776 15206
rect 17468 15195 17776 15204
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17236 14742 17356 14770
rect 16948 14554 17000 14560
rect 17052 14572 17172 14600
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16684 12850 16712 14418
rect 16960 13870 16988 14554
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17052 13734 17080 14572
rect 17328 14464 17356 14742
rect 17512 14618 17540 14962
rect 17880 14906 17908 19994
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17972 18222 18000 19926
rect 18156 19854 18184 21714
rect 18708 19854 18736 21714
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18064 17338 18092 17546
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18156 15978 18184 16934
rect 18248 16538 18276 19654
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18834 18460 19110
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18524 18358 18552 18838
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18524 17882 18552 18294
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18248 16510 18368 16538
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18248 16250 18276 16390
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18236 14952 18288 14958
rect 17880 14878 18000 14906
rect 18236 14894 18288 14900
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17144 14436 17356 14464
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16808 13628 17116 13637
rect 16808 13626 16814 13628
rect 16870 13626 16894 13628
rect 16950 13626 16974 13628
rect 17030 13626 17054 13628
rect 17110 13626 17116 13628
rect 16870 13574 16872 13626
rect 17052 13574 17054 13626
rect 16808 13572 16814 13574
rect 16870 13572 16894 13574
rect 16950 13572 16974 13574
rect 17030 13572 17054 13574
rect 17110 13572 17116 13574
rect 16808 13563 17116 13572
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16684 12306 16712 12650
rect 16808 12540 17116 12549
rect 16808 12538 16814 12540
rect 16870 12538 16894 12540
rect 16950 12538 16974 12540
rect 17030 12538 17054 12540
rect 17110 12538 17116 12540
rect 16870 12486 16872 12538
rect 17052 12486 17054 12538
rect 16808 12484 16814 12486
rect 16870 12484 16894 12486
rect 16950 12484 16974 12486
rect 17030 12484 17054 12486
rect 17110 12484 17116 12486
rect 16808 12475 17116 12484
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16868 11898 16896 12038
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16808 11452 17116 11461
rect 16808 11450 16814 11452
rect 16870 11450 16894 11452
rect 16950 11450 16974 11452
rect 17030 11450 17054 11452
rect 17110 11450 17116 11452
rect 16870 11398 16872 11450
rect 17052 11398 17054 11450
rect 16808 11396 16814 11398
rect 16870 11396 16894 11398
rect 16950 11396 16974 11398
rect 17030 11396 17054 11398
rect 17110 11396 17116 11398
rect 16808 11387 17116 11396
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16500 10062 16528 10610
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 10266 16620 10474
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9722 16528 9862
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16224 9178 16252 9454
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15396 6866 15424 7278
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15488 6798 15516 7686
rect 15580 6798 15608 8366
rect 15856 8090 15884 8910
rect 16408 8498 16436 8910
rect 16500 8566 16528 9658
rect 16684 9586 16712 10542
rect 16808 10364 17116 10373
rect 16808 10362 16814 10364
rect 16870 10362 16894 10364
rect 16950 10362 16974 10364
rect 17030 10362 17054 10364
rect 17110 10362 17116 10364
rect 16870 10310 16872 10362
rect 17052 10310 17054 10362
rect 16808 10308 16814 10310
rect 16870 10308 16894 10310
rect 16950 10308 16974 10310
rect 17030 10308 17054 10310
rect 17110 10308 17116 10310
rect 16808 10299 17116 10308
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 16408 7886 16436 8434
rect 16592 8362 16620 8978
rect 16684 8498 16712 9522
rect 16808 9276 17116 9285
rect 16808 9274 16814 9276
rect 16870 9274 16894 9276
rect 16950 9274 16974 9276
rect 17030 9274 17054 9276
rect 17110 9274 17116 9276
rect 16870 9222 16872 9274
rect 17052 9222 17054 9274
rect 16808 9220 16814 9222
rect 16870 9220 16894 9222
rect 16950 9220 16974 9222
rect 17030 9220 17054 9222
rect 17110 9220 17116 9222
rect 16808 9211 17116 9220
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16808 8188 17116 8197
rect 16808 8186 16814 8188
rect 16870 8186 16894 8188
rect 16950 8186 16974 8188
rect 17030 8186 17054 8188
rect 17110 8186 17116 8188
rect 16870 8134 16872 8186
rect 17052 8134 17054 8186
rect 16808 8132 16814 8134
rect 16870 8132 16894 8134
rect 16950 8132 16974 8134
rect 17030 8132 17054 8134
rect 17110 8132 17116 8134
rect 16808 8123 17116 8132
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 17144 7546 17172 14436
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13410 17264 13670
rect 17328 13530 17356 14282
rect 17468 14172 17776 14181
rect 17468 14170 17474 14172
rect 17530 14170 17554 14172
rect 17610 14170 17634 14172
rect 17690 14170 17714 14172
rect 17770 14170 17776 14172
rect 17530 14118 17532 14170
rect 17712 14118 17714 14170
rect 17468 14116 17474 14118
rect 17530 14116 17554 14118
rect 17610 14116 17634 14118
rect 17690 14116 17714 14118
rect 17770 14116 17776 14118
rect 17468 14107 17776 14116
rect 17880 14006 17908 14758
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17236 13382 17356 13410
rect 17880 13394 17908 13942
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17236 11694 17264 12242
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17328 8090 17356 13382
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17972 13274 18000 14878
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 14074 18092 14214
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18248 13938 18276 14894
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 17880 13246 18000 13274
rect 17468 13084 17776 13093
rect 17468 13082 17474 13084
rect 17530 13082 17554 13084
rect 17610 13082 17634 13084
rect 17690 13082 17714 13084
rect 17770 13082 17776 13084
rect 17530 13030 17532 13082
rect 17712 13030 17714 13082
rect 17468 13028 17474 13030
rect 17530 13028 17554 13030
rect 17610 13028 17634 13030
rect 17690 13028 17714 13030
rect 17770 13028 17776 13030
rect 17468 13019 17776 13028
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17420 12374 17448 12718
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17468 11996 17776 12005
rect 17468 11994 17474 11996
rect 17530 11994 17554 11996
rect 17610 11994 17634 11996
rect 17690 11994 17714 11996
rect 17770 11994 17776 11996
rect 17530 11942 17532 11994
rect 17712 11942 17714 11994
rect 17468 11940 17474 11942
rect 17530 11940 17554 11942
rect 17610 11940 17634 11942
rect 17690 11940 17714 11942
rect 17770 11940 17776 11942
rect 17468 11931 17776 11940
rect 17468 10908 17776 10917
rect 17468 10906 17474 10908
rect 17530 10906 17554 10908
rect 17610 10906 17634 10908
rect 17690 10906 17714 10908
rect 17770 10906 17776 10908
rect 17530 10854 17532 10906
rect 17712 10854 17714 10906
rect 17468 10852 17474 10854
rect 17530 10852 17554 10854
rect 17610 10852 17634 10854
rect 17690 10852 17714 10854
rect 17770 10852 17776 10854
rect 17468 10843 17776 10852
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10062 17540 10406
rect 17696 10266 17724 10678
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17468 9820 17776 9829
rect 17468 9818 17474 9820
rect 17530 9818 17554 9820
rect 17610 9818 17634 9820
rect 17690 9818 17714 9820
rect 17770 9818 17776 9820
rect 17530 9766 17532 9818
rect 17712 9766 17714 9818
rect 17468 9764 17474 9766
rect 17530 9764 17554 9766
rect 17610 9764 17634 9766
rect 17690 9764 17714 9766
rect 17770 9764 17776 9766
rect 17468 9755 17776 9764
rect 17880 8974 17908 13246
rect 18248 12986 18276 13874
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12238 18092 12582
rect 18340 12434 18368 16510
rect 18524 16114 18552 16594
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18524 14074 18552 14350
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18432 12442 18460 12854
rect 18156 12406 18368 12434
rect 18420 12436 18472 12442
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 9926 18000 12038
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17972 9518 18000 9862
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17972 8786 18000 9454
rect 17880 8758 18000 8786
rect 17468 8732 17776 8741
rect 17468 8730 17474 8732
rect 17530 8730 17554 8732
rect 17610 8730 17634 8732
rect 17690 8730 17714 8732
rect 17770 8730 17776 8732
rect 17530 8678 17532 8730
rect 17712 8678 17714 8730
rect 17468 8676 17474 8678
rect 17530 8676 17554 8678
rect 17610 8676 17634 8678
rect 17690 8676 17714 8678
rect 17770 8676 17776 8678
rect 17468 8667 17776 8676
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17420 8090 17448 8502
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17604 8090 17632 8230
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17880 7818 17908 8758
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17468 7644 17776 7653
rect 17468 7642 17474 7644
rect 17530 7642 17554 7644
rect 17610 7642 17634 7644
rect 17690 7642 17714 7644
rect 17770 7642 17776 7644
rect 17530 7590 17532 7642
rect 17712 7590 17714 7642
rect 17468 7588 17474 7590
rect 17530 7588 17554 7590
rect 17610 7588 17634 7590
rect 17690 7588 17714 7590
rect 17770 7588 17776 7590
rect 17468 7579 17776 7588
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14660 5370 14688 6394
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13280 4826 13308 5238
rect 14936 5166 14964 6598
rect 15580 6390 15608 6598
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15856 6322 15884 6598
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15948 6118 15976 6666
rect 16592 6662 16620 7278
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 16040 5846 16068 6598
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 16224 5710 16252 6122
rect 16316 5778 16344 6258
rect 16684 5914 16712 7142
rect 16808 7100 17116 7109
rect 16808 7098 16814 7100
rect 16870 7098 16894 7100
rect 16950 7098 16974 7100
rect 17030 7098 17054 7100
rect 17110 7098 17116 7100
rect 16870 7046 16872 7098
rect 17052 7046 17054 7098
rect 16808 7044 16814 7046
rect 16870 7044 16894 7046
rect 16950 7044 16974 7046
rect 17030 7044 17054 7046
rect 17110 7044 17116 7046
rect 16808 7035 17116 7044
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16776 6390 16804 6734
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16868 6186 16896 6802
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 6390 17080 6598
rect 17468 6556 17776 6565
rect 17468 6554 17474 6556
rect 17530 6554 17554 6556
rect 17610 6554 17634 6556
rect 17690 6554 17714 6556
rect 17770 6554 17776 6556
rect 17530 6502 17532 6554
rect 17712 6502 17714 6554
rect 17468 6500 17474 6502
rect 17530 6500 17554 6502
rect 17610 6500 17634 6502
rect 17690 6500 17714 6502
rect 17770 6500 17776 6502
rect 17468 6491 17776 6500
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16808 6012 17116 6021
rect 16808 6010 16814 6012
rect 16870 6010 16894 6012
rect 16950 6010 16974 6012
rect 17030 6010 17054 6012
rect 17110 6010 17116 6012
rect 16870 5958 16872 6010
rect 17052 5958 17054 6010
rect 16808 5956 16814 5958
rect 16870 5956 16894 5958
rect 16950 5956 16974 5958
rect 17030 5956 17054 5958
rect 17110 5956 17116 5958
rect 16808 5947 17116 5956
rect 17420 5914 17448 6326
rect 17880 6118 17908 7754
rect 18156 6254 18184 12406
rect 18708 12434 18736 19654
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18892 14618 18920 15982
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18420 12378 18472 12384
rect 18616 12406 18736 12434
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18340 10810 18368 11086
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18340 10062 18368 10746
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 7954 18460 8230
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18524 7546 18552 8570
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18616 7206 18644 12406
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10674 18920 10950
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18708 10130 18736 10610
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18708 9722 18736 10066
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18800 7410 18828 7890
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18800 6458 18828 7346
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16316 5370 16344 5714
rect 17880 5710 17908 6054
rect 18432 5914 18460 6326
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17468 5468 17776 5477
rect 17468 5466 17474 5468
rect 17530 5466 17554 5468
rect 17610 5466 17634 5468
rect 17690 5466 17714 5468
rect 17770 5466 17776 5468
rect 17530 5414 17532 5466
rect 17712 5414 17714 5466
rect 17468 5412 17474 5414
rect 17530 5412 17554 5414
rect 17610 5412 17634 5414
rect 17690 5412 17714 5414
rect 17770 5412 17776 5414
rect 17468 5403 17776 5412
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15120 4826 15148 5238
rect 16808 4924 17116 4933
rect 16808 4922 16814 4924
rect 16870 4922 16894 4924
rect 16950 4922 16974 4924
rect 17030 4922 17054 4924
rect 17110 4922 17116 4924
rect 16870 4870 16872 4922
rect 17052 4870 17054 4922
rect 16808 4868 16814 4870
rect 16870 4868 16894 4870
rect 16950 4868 16974 4870
rect 17030 4868 17054 4870
rect 17110 4868 17116 4870
rect 16808 4859 17116 4868
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2792 4282 2820 4490
rect 3875 4380 4183 4389
rect 3875 4378 3881 4380
rect 3937 4378 3961 4380
rect 4017 4378 4041 4380
rect 4097 4378 4121 4380
rect 4177 4378 4183 4380
rect 3937 4326 3939 4378
rect 4119 4326 4121 4378
rect 3875 4324 3881 4326
rect 3937 4324 3961 4326
rect 4017 4324 4041 4326
rect 4097 4324 4121 4326
rect 4177 4324 4183 4326
rect 3875 4315 4183 4324
rect 8406 4380 8714 4389
rect 8406 4378 8412 4380
rect 8468 4378 8492 4380
rect 8548 4378 8572 4380
rect 8628 4378 8652 4380
rect 8708 4378 8714 4380
rect 8468 4326 8470 4378
rect 8650 4326 8652 4378
rect 8406 4324 8412 4326
rect 8468 4324 8492 4326
rect 8548 4324 8572 4326
rect 8628 4324 8652 4326
rect 8708 4324 8714 4326
rect 8406 4315 8714 4324
rect 12937 4380 13245 4389
rect 12937 4378 12943 4380
rect 12999 4378 13023 4380
rect 13079 4378 13103 4380
rect 13159 4378 13183 4380
rect 13239 4378 13245 4380
rect 12999 4326 13001 4378
rect 13181 4326 13183 4378
rect 12937 4324 12943 4326
rect 12999 4324 13023 4326
rect 13079 4324 13103 4326
rect 13159 4324 13183 4326
rect 13239 4324 13245 4326
rect 12937 4315 13245 4324
rect 14936 4282 14964 4558
rect 17468 4380 17776 4389
rect 17468 4378 17474 4380
rect 17530 4378 17554 4380
rect 17610 4378 17634 4380
rect 17690 4378 17714 4380
rect 17770 4378 17776 4380
rect 17530 4326 17532 4378
rect 17712 4326 17714 4378
rect 17468 4324 17474 4326
rect 17530 4324 17554 4326
rect 17610 4324 17634 4326
rect 17690 4324 17714 4326
rect 17770 4324 17776 4326
rect 17468 4315 17776 4324
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 3215 3836 3523 3845
rect 3215 3834 3221 3836
rect 3277 3834 3301 3836
rect 3357 3834 3381 3836
rect 3437 3834 3461 3836
rect 3517 3834 3523 3836
rect 3277 3782 3279 3834
rect 3459 3782 3461 3834
rect 3215 3780 3221 3782
rect 3277 3780 3301 3782
rect 3357 3780 3381 3782
rect 3437 3780 3461 3782
rect 3517 3780 3523 3782
rect 3215 3771 3523 3780
rect 7746 3836 8054 3845
rect 7746 3834 7752 3836
rect 7808 3834 7832 3836
rect 7888 3834 7912 3836
rect 7968 3834 7992 3836
rect 8048 3834 8054 3836
rect 7808 3782 7810 3834
rect 7990 3782 7992 3834
rect 7746 3780 7752 3782
rect 7808 3780 7832 3782
rect 7888 3780 7912 3782
rect 7968 3780 7992 3782
rect 8048 3780 8054 3782
rect 7746 3771 8054 3780
rect 12277 3836 12585 3845
rect 12277 3834 12283 3836
rect 12339 3834 12363 3836
rect 12419 3834 12443 3836
rect 12499 3834 12523 3836
rect 12579 3834 12585 3836
rect 12339 3782 12341 3834
rect 12521 3782 12523 3834
rect 12277 3780 12283 3782
rect 12339 3780 12363 3782
rect 12419 3780 12443 3782
rect 12499 3780 12523 3782
rect 12579 3780 12585 3782
rect 12277 3771 12585 3780
rect 3875 3292 4183 3301
rect 3875 3290 3881 3292
rect 3937 3290 3961 3292
rect 4017 3290 4041 3292
rect 4097 3290 4121 3292
rect 4177 3290 4183 3292
rect 3937 3238 3939 3290
rect 4119 3238 4121 3290
rect 3875 3236 3881 3238
rect 3937 3236 3961 3238
rect 4017 3236 4041 3238
rect 4097 3236 4121 3238
rect 4177 3236 4183 3238
rect 3875 3227 4183 3236
rect 8406 3292 8714 3301
rect 8406 3290 8412 3292
rect 8468 3290 8492 3292
rect 8548 3290 8572 3292
rect 8628 3290 8652 3292
rect 8708 3290 8714 3292
rect 8468 3238 8470 3290
rect 8650 3238 8652 3290
rect 8406 3236 8412 3238
rect 8468 3236 8492 3238
rect 8548 3236 8572 3238
rect 8628 3236 8652 3238
rect 8708 3236 8714 3238
rect 8406 3227 8714 3236
rect 12937 3292 13245 3301
rect 12937 3290 12943 3292
rect 12999 3290 13023 3292
rect 13079 3290 13103 3292
rect 13159 3290 13183 3292
rect 13239 3290 13245 3292
rect 12999 3238 13001 3290
rect 13181 3238 13183 3290
rect 12937 3236 12943 3238
rect 12999 3236 13023 3238
rect 13079 3236 13103 3238
rect 13159 3236 13183 3238
rect 13239 3236 13245 3238
rect 12937 3227 13245 3236
rect 3215 2748 3523 2757
rect 3215 2746 3221 2748
rect 3277 2746 3301 2748
rect 3357 2746 3381 2748
rect 3437 2746 3461 2748
rect 3517 2746 3523 2748
rect 3277 2694 3279 2746
rect 3459 2694 3461 2746
rect 3215 2692 3221 2694
rect 3277 2692 3301 2694
rect 3357 2692 3381 2694
rect 3437 2692 3461 2694
rect 3517 2692 3523 2694
rect 3215 2683 3523 2692
rect 7746 2748 8054 2757
rect 7746 2746 7752 2748
rect 7808 2746 7832 2748
rect 7888 2746 7912 2748
rect 7968 2746 7992 2748
rect 8048 2746 8054 2748
rect 7808 2694 7810 2746
rect 7990 2694 7992 2746
rect 7746 2692 7752 2694
rect 7808 2692 7832 2694
rect 7888 2692 7912 2694
rect 7968 2692 7992 2694
rect 8048 2692 8054 2694
rect 7746 2683 8054 2692
rect 12277 2748 12585 2757
rect 12277 2746 12283 2748
rect 12339 2746 12363 2748
rect 12419 2746 12443 2748
rect 12499 2746 12523 2748
rect 12579 2746 12585 2748
rect 12339 2694 12341 2746
rect 12521 2694 12523 2746
rect 12277 2692 12283 2694
rect 12339 2692 12363 2694
rect 12419 2692 12443 2694
rect 12499 2692 12523 2694
rect 12579 2692 12585 2694
rect 12277 2683 12585 2692
rect 15304 2650 15332 4150
rect 16808 3836 17116 3845
rect 16808 3834 16814 3836
rect 16870 3834 16894 3836
rect 16950 3834 16974 3836
rect 17030 3834 17054 3836
rect 17110 3834 17116 3836
rect 16870 3782 16872 3834
rect 17052 3782 17054 3834
rect 16808 3780 16814 3782
rect 16870 3780 16894 3782
rect 16950 3780 16974 3782
rect 17030 3780 17054 3782
rect 17110 3780 17116 3782
rect 16808 3771 17116 3780
rect 17468 3292 17776 3301
rect 17468 3290 17474 3292
rect 17530 3290 17554 3292
rect 17610 3290 17634 3292
rect 17690 3290 17714 3292
rect 17770 3290 17776 3292
rect 17530 3238 17532 3290
rect 17712 3238 17714 3290
rect 17468 3236 17474 3238
rect 17530 3236 17554 3238
rect 17610 3236 17634 3238
rect 17690 3236 17714 3238
rect 17770 3236 17776 3238
rect 17468 3227 17776 3236
rect 16808 2748 17116 2757
rect 16808 2746 16814 2748
rect 16870 2746 16894 2748
rect 16950 2746 16974 2748
rect 17030 2746 17054 2748
rect 17110 2746 17116 2748
rect 16870 2694 16872 2746
rect 17052 2694 17054 2746
rect 16808 2692 16814 2694
rect 16870 2692 16894 2694
rect 16950 2692 16974 2694
rect 17030 2692 17054 2694
rect 17110 2692 17116 2694
rect 16808 2683 17116 2692
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 3875 2204 4183 2213
rect 3875 2202 3881 2204
rect 3937 2202 3961 2204
rect 4017 2202 4041 2204
rect 4097 2202 4121 2204
rect 4177 2202 4183 2204
rect 3937 2150 3939 2202
rect 4119 2150 4121 2202
rect 3875 2148 3881 2150
rect 3937 2148 3961 2150
rect 4017 2148 4041 2150
rect 4097 2148 4121 2150
rect 4177 2148 4183 2150
rect 3875 2139 4183 2148
rect 8406 2204 8714 2213
rect 8406 2202 8412 2204
rect 8468 2202 8492 2204
rect 8548 2202 8572 2204
rect 8628 2202 8652 2204
rect 8708 2202 8714 2204
rect 8468 2150 8470 2202
rect 8650 2150 8652 2202
rect 8406 2148 8412 2150
rect 8468 2148 8492 2150
rect 8548 2148 8572 2150
rect 8628 2148 8652 2150
rect 8708 2148 8714 2150
rect 8406 2139 8714 2148
rect 12937 2204 13245 2213
rect 12937 2202 12943 2204
rect 12999 2202 13023 2204
rect 13079 2202 13103 2204
rect 13159 2202 13183 2204
rect 13239 2202 13245 2204
rect 12999 2150 13001 2202
rect 13181 2150 13183 2202
rect 12937 2148 12943 2150
rect 12999 2148 13023 2150
rect 13079 2148 13103 2150
rect 13159 2148 13183 2150
rect 13239 2148 13245 2150
rect 12937 2139 13245 2148
rect 15304 1306 15332 2382
rect 17468 2204 17776 2213
rect 17468 2202 17474 2204
rect 17530 2202 17554 2204
rect 17610 2202 17634 2204
rect 17690 2202 17714 2204
rect 17770 2202 17776 2204
rect 17530 2150 17532 2202
rect 17712 2150 17714 2202
rect 17468 2148 17474 2150
rect 17530 2148 17554 2150
rect 17610 2148 17634 2150
rect 17690 2148 17714 2150
rect 17770 2148 17776 2150
rect 17468 2139 17776 2148
rect 15212 1278 15332 1306
rect 15212 800 15240 1278
rect 15198 0 15254 800
<< via2 >>
rect 938 16632 994 16688
rect 3221 20154 3277 20156
rect 3301 20154 3357 20156
rect 3381 20154 3437 20156
rect 3461 20154 3517 20156
rect 3221 20102 3267 20154
rect 3267 20102 3277 20154
rect 3301 20102 3331 20154
rect 3331 20102 3343 20154
rect 3343 20102 3357 20154
rect 3381 20102 3395 20154
rect 3395 20102 3407 20154
rect 3407 20102 3437 20154
rect 3461 20102 3471 20154
rect 3471 20102 3517 20154
rect 3221 20100 3277 20102
rect 3301 20100 3357 20102
rect 3381 20100 3437 20102
rect 3461 20100 3517 20102
rect 7752 20154 7808 20156
rect 7832 20154 7888 20156
rect 7912 20154 7968 20156
rect 7992 20154 8048 20156
rect 7752 20102 7798 20154
rect 7798 20102 7808 20154
rect 7832 20102 7862 20154
rect 7862 20102 7874 20154
rect 7874 20102 7888 20154
rect 7912 20102 7926 20154
rect 7926 20102 7938 20154
rect 7938 20102 7968 20154
rect 7992 20102 8002 20154
rect 8002 20102 8048 20154
rect 7752 20100 7808 20102
rect 7832 20100 7888 20102
rect 7912 20100 7968 20102
rect 7992 20100 8048 20102
rect 3881 19610 3937 19612
rect 3961 19610 4017 19612
rect 4041 19610 4097 19612
rect 4121 19610 4177 19612
rect 3881 19558 3927 19610
rect 3927 19558 3937 19610
rect 3961 19558 3991 19610
rect 3991 19558 4003 19610
rect 4003 19558 4017 19610
rect 4041 19558 4055 19610
rect 4055 19558 4067 19610
rect 4067 19558 4097 19610
rect 4121 19558 4131 19610
rect 4131 19558 4177 19610
rect 3881 19556 3937 19558
rect 3961 19556 4017 19558
rect 4041 19556 4097 19558
rect 4121 19556 4177 19558
rect 3221 19066 3277 19068
rect 3301 19066 3357 19068
rect 3381 19066 3437 19068
rect 3461 19066 3517 19068
rect 3221 19014 3267 19066
rect 3267 19014 3277 19066
rect 3301 19014 3331 19066
rect 3331 19014 3343 19066
rect 3343 19014 3357 19066
rect 3381 19014 3395 19066
rect 3395 19014 3407 19066
rect 3407 19014 3437 19066
rect 3461 19014 3471 19066
rect 3471 19014 3517 19066
rect 3221 19012 3277 19014
rect 3301 19012 3357 19014
rect 3381 19012 3437 19014
rect 3461 19012 3517 19014
rect 3881 18522 3937 18524
rect 3961 18522 4017 18524
rect 4041 18522 4097 18524
rect 4121 18522 4177 18524
rect 3881 18470 3927 18522
rect 3927 18470 3937 18522
rect 3961 18470 3991 18522
rect 3991 18470 4003 18522
rect 4003 18470 4017 18522
rect 4041 18470 4055 18522
rect 4055 18470 4067 18522
rect 4067 18470 4097 18522
rect 4121 18470 4131 18522
rect 4131 18470 4177 18522
rect 3881 18468 3937 18470
rect 3961 18468 4017 18470
rect 4041 18468 4097 18470
rect 4121 18468 4177 18470
rect 3221 17978 3277 17980
rect 3301 17978 3357 17980
rect 3381 17978 3437 17980
rect 3461 17978 3517 17980
rect 3221 17926 3267 17978
rect 3267 17926 3277 17978
rect 3301 17926 3331 17978
rect 3331 17926 3343 17978
rect 3343 17926 3357 17978
rect 3381 17926 3395 17978
rect 3395 17926 3407 17978
rect 3407 17926 3437 17978
rect 3461 17926 3471 17978
rect 3471 17926 3517 17978
rect 3221 17924 3277 17926
rect 3301 17924 3357 17926
rect 3381 17924 3437 17926
rect 3461 17924 3517 17926
rect 3221 16890 3277 16892
rect 3301 16890 3357 16892
rect 3381 16890 3437 16892
rect 3461 16890 3517 16892
rect 3221 16838 3267 16890
rect 3267 16838 3277 16890
rect 3301 16838 3331 16890
rect 3331 16838 3343 16890
rect 3343 16838 3357 16890
rect 3381 16838 3395 16890
rect 3395 16838 3407 16890
rect 3407 16838 3437 16890
rect 3461 16838 3471 16890
rect 3471 16838 3517 16890
rect 3221 16836 3277 16838
rect 3301 16836 3357 16838
rect 3381 16836 3437 16838
rect 3461 16836 3517 16838
rect 2686 12844 2742 12880
rect 2686 12824 2688 12844
rect 2688 12824 2740 12844
rect 2740 12824 2742 12844
rect 3221 15802 3277 15804
rect 3301 15802 3357 15804
rect 3381 15802 3437 15804
rect 3461 15802 3517 15804
rect 3221 15750 3267 15802
rect 3267 15750 3277 15802
rect 3301 15750 3331 15802
rect 3331 15750 3343 15802
rect 3343 15750 3357 15802
rect 3381 15750 3395 15802
rect 3395 15750 3407 15802
rect 3407 15750 3437 15802
rect 3461 15750 3471 15802
rect 3471 15750 3517 15802
rect 3221 15748 3277 15750
rect 3301 15748 3357 15750
rect 3381 15748 3437 15750
rect 3461 15748 3517 15750
rect 3221 14714 3277 14716
rect 3301 14714 3357 14716
rect 3381 14714 3437 14716
rect 3461 14714 3517 14716
rect 3221 14662 3267 14714
rect 3267 14662 3277 14714
rect 3301 14662 3331 14714
rect 3331 14662 3343 14714
rect 3343 14662 3357 14714
rect 3381 14662 3395 14714
rect 3395 14662 3407 14714
rect 3407 14662 3437 14714
rect 3461 14662 3471 14714
rect 3471 14662 3517 14714
rect 3221 14660 3277 14662
rect 3301 14660 3357 14662
rect 3381 14660 3437 14662
rect 3461 14660 3517 14662
rect 3221 13626 3277 13628
rect 3301 13626 3357 13628
rect 3381 13626 3437 13628
rect 3461 13626 3517 13628
rect 3221 13574 3267 13626
rect 3267 13574 3277 13626
rect 3301 13574 3331 13626
rect 3331 13574 3343 13626
rect 3343 13574 3357 13626
rect 3381 13574 3395 13626
rect 3395 13574 3407 13626
rect 3407 13574 3437 13626
rect 3461 13574 3471 13626
rect 3471 13574 3517 13626
rect 3221 13572 3277 13574
rect 3301 13572 3357 13574
rect 3381 13572 3437 13574
rect 3461 13572 3517 13574
rect 3881 17434 3937 17436
rect 3961 17434 4017 17436
rect 4041 17434 4097 17436
rect 4121 17434 4177 17436
rect 3881 17382 3927 17434
rect 3927 17382 3937 17434
rect 3961 17382 3991 17434
rect 3991 17382 4003 17434
rect 4003 17382 4017 17434
rect 4041 17382 4055 17434
rect 4055 17382 4067 17434
rect 4067 17382 4097 17434
rect 4121 17382 4131 17434
rect 4131 17382 4177 17434
rect 3881 17380 3937 17382
rect 3961 17380 4017 17382
rect 4041 17380 4097 17382
rect 4121 17380 4177 17382
rect 3881 16346 3937 16348
rect 3961 16346 4017 16348
rect 4041 16346 4097 16348
rect 4121 16346 4177 16348
rect 3881 16294 3927 16346
rect 3927 16294 3937 16346
rect 3961 16294 3991 16346
rect 3991 16294 4003 16346
rect 4003 16294 4017 16346
rect 4041 16294 4055 16346
rect 4055 16294 4067 16346
rect 4067 16294 4097 16346
rect 4121 16294 4131 16346
rect 4131 16294 4177 16346
rect 3881 16292 3937 16294
rect 3961 16292 4017 16294
rect 4041 16292 4097 16294
rect 4121 16292 4177 16294
rect 3881 15258 3937 15260
rect 3961 15258 4017 15260
rect 4041 15258 4097 15260
rect 4121 15258 4177 15260
rect 3881 15206 3927 15258
rect 3927 15206 3937 15258
rect 3961 15206 3991 15258
rect 3991 15206 4003 15258
rect 4003 15206 4017 15258
rect 4041 15206 4055 15258
rect 4055 15206 4067 15258
rect 4067 15206 4097 15258
rect 4121 15206 4131 15258
rect 4131 15206 4177 15258
rect 3881 15204 3937 15206
rect 3961 15204 4017 15206
rect 4041 15204 4097 15206
rect 4121 15204 4177 15206
rect 3881 14170 3937 14172
rect 3961 14170 4017 14172
rect 4041 14170 4097 14172
rect 4121 14170 4177 14172
rect 3881 14118 3927 14170
rect 3927 14118 3937 14170
rect 3961 14118 3991 14170
rect 3991 14118 4003 14170
rect 4003 14118 4017 14170
rect 4041 14118 4055 14170
rect 4055 14118 4067 14170
rect 4067 14118 4097 14170
rect 4121 14118 4131 14170
rect 4131 14118 4177 14170
rect 3881 14116 3937 14118
rect 3961 14116 4017 14118
rect 4041 14116 4097 14118
rect 4121 14116 4177 14118
rect 3881 13082 3937 13084
rect 3961 13082 4017 13084
rect 4041 13082 4097 13084
rect 4121 13082 4177 13084
rect 3881 13030 3927 13082
rect 3927 13030 3937 13082
rect 3961 13030 3991 13082
rect 3991 13030 4003 13082
rect 4003 13030 4017 13082
rect 4041 13030 4055 13082
rect 4055 13030 4067 13082
rect 4067 13030 4097 13082
rect 4121 13030 4131 13082
rect 4131 13030 4177 13082
rect 3881 13028 3937 13030
rect 3961 13028 4017 13030
rect 4041 13028 4097 13030
rect 4121 13028 4177 13030
rect 3221 12538 3277 12540
rect 3301 12538 3357 12540
rect 3381 12538 3437 12540
rect 3461 12538 3517 12540
rect 3221 12486 3267 12538
rect 3267 12486 3277 12538
rect 3301 12486 3331 12538
rect 3331 12486 3343 12538
rect 3343 12486 3357 12538
rect 3381 12486 3395 12538
rect 3395 12486 3407 12538
rect 3407 12486 3437 12538
rect 3461 12486 3471 12538
rect 3471 12486 3517 12538
rect 3221 12484 3277 12486
rect 3301 12484 3357 12486
rect 3381 12484 3437 12486
rect 3461 12484 3517 12486
rect 3221 11450 3277 11452
rect 3301 11450 3357 11452
rect 3381 11450 3437 11452
rect 3461 11450 3517 11452
rect 3221 11398 3267 11450
rect 3267 11398 3277 11450
rect 3301 11398 3331 11450
rect 3331 11398 3343 11450
rect 3343 11398 3357 11450
rect 3381 11398 3395 11450
rect 3395 11398 3407 11450
rect 3407 11398 3437 11450
rect 3461 11398 3471 11450
rect 3471 11398 3517 11450
rect 3221 11396 3277 11398
rect 3301 11396 3357 11398
rect 3381 11396 3437 11398
rect 3461 11396 3517 11398
rect 3221 10362 3277 10364
rect 3301 10362 3357 10364
rect 3381 10362 3437 10364
rect 3461 10362 3517 10364
rect 3221 10310 3267 10362
rect 3267 10310 3277 10362
rect 3301 10310 3331 10362
rect 3331 10310 3343 10362
rect 3343 10310 3357 10362
rect 3381 10310 3395 10362
rect 3395 10310 3407 10362
rect 3407 10310 3437 10362
rect 3461 10310 3471 10362
rect 3471 10310 3517 10362
rect 3221 10308 3277 10310
rect 3301 10308 3357 10310
rect 3381 10308 3437 10310
rect 3461 10308 3517 10310
rect 3221 9274 3277 9276
rect 3301 9274 3357 9276
rect 3381 9274 3437 9276
rect 3461 9274 3517 9276
rect 3221 9222 3267 9274
rect 3267 9222 3277 9274
rect 3301 9222 3331 9274
rect 3331 9222 3343 9274
rect 3343 9222 3357 9274
rect 3381 9222 3395 9274
rect 3395 9222 3407 9274
rect 3407 9222 3437 9274
rect 3461 9222 3471 9274
rect 3471 9222 3517 9274
rect 3221 9220 3277 9222
rect 3301 9220 3357 9222
rect 3381 9220 3437 9222
rect 3461 9220 3517 9222
rect 3881 11994 3937 11996
rect 3961 11994 4017 11996
rect 4041 11994 4097 11996
rect 4121 11994 4177 11996
rect 3881 11942 3927 11994
rect 3927 11942 3937 11994
rect 3961 11942 3991 11994
rect 3991 11942 4003 11994
rect 4003 11942 4017 11994
rect 4041 11942 4055 11994
rect 4055 11942 4067 11994
rect 4067 11942 4097 11994
rect 4121 11942 4131 11994
rect 4131 11942 4177 11994
rect 3881 11940 3937 11942
rect 3961 11940 4017 11942
rect 4041 11940 4097 11942
rect 4121 11940 4177 11942
rect 3881 10906 3937 10908
rect 3961 10906 4017 10908
rect 4041 10906 4097 10908
rect 4121 10906 4177 10908
rect 3881 10854 3927 10906
rect 3927 10854 3937 10906
rect 3961 10854 3991 10906
rect 3991 10854 4003 10906
rect 4003 10854 4017 10906
rect 4041 10854 4055 10906
rect 4055 10854 4067 10906
rect 4067 10854 4097 10906
rect 4121 10854 4131 10906
rect 4131 10854 4177 10906
rect 3881 10852 3937 10854
rect 3961 10852 4017 10854
rect 4041 10852 4097 10854
rect 4121 10852 4177 10854
rect 3881 9818 3937 9820
rect 3961 9818 4017 9820
rect 4041 9818 4097 9820
rect 4121 9818 4177 9820
rect 3881 9766 3927 9818
rect 3927 9766 3937 9818
rect 3961 9766 3991 9818
rect 3991 9766 4003 9818
rect 4003 9766 4017 9818
rect 4041 9766 4055 9818
rect 4055 9766 4067 9818
rect 4067 9766 4097 9818
rect 4121 9766 4131 9818
rect 4131 9766 4177 9818
rect 3881 9764 3937 9766
rect 3961 9764 4017 9766
rect 4041 9764 4097 9766
rect 4121 9764 4177 9766
rect 3881 8730 3937 8732
rect 3961 8730 4017 8732
rect 4041 8730 4097 8732
rect 4121 8730 4177 8732
rect 3881 8678 3927 8730
rect 3927 8678 3937 8730
rect 3961 8678 3991 8730
rect 3991 8678 4003 8730
rect 4003 8678 4017 8730
rect 4041 8678 4055 8730
rect 4055 8678 4067 8730
rect 4067 8678 4097 8730
rect 4121 8678 4131 8730
rect 4131 8678 4177 8730
rect 3881 8676 3937 8678
rect 3961 8676 4017 8678
rect 4041 8676 4097 8678
rect 4121 8676 4177 8678
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 4158 8200 4214 8256
rect 3221 8186 3277 8188
rect 3301 8186 3357 8188
rect 3381 8186 3437 8188
rect 3461 8186 3517 8188
rect 3221 8134 3267 8186
rect 3267 8134 3277 8186
rect 3301 8134 3331 8186
rect 3331 8134 3343 8186
rect 3343 8134 3357 8186
rect 3381 8134 3395 8186
rect 3395 8134 3407 8186
rect 3407 8134 3437 8186
rect 3461 8134 3471 8186
rect 3471 8134 3517 8186
rect 3221 8132 3277 8134
rect 3301 8132 3357 8134
rect 3381 8132 3437 8134
rect 3461 8132 3517 8134
rect 3881 7642 3937 7644
rect 3961 7642 4017 7644
rect 4041 7642 4097 7644
rect 4121 7642 4177 7644
rect 3881 7590 3927 7642
rect 3927 7590 3937 7642
rect 3961 7590 3991 7642
rect 3991 7590 4003 7642
rect 4003 7590 4017 7642
rect 4041 7590 4055 7642
rect 4055 7590 4067 7642
rect 4067 7590 4097 7642
rect 4121 7590 4131 7642
rect 4131 7590 4177 7642
rect 3881 7588 3937 7590
rect 3961 7588 4017 7590
rect 4041 7588 4097 7590
rect 4121 7588 4177 7590
rect 8412 19610 8468 19612
rect 8492 19610 8548 19612
rect 8572 19610 8628 19612
rect 8652 19610 8708 19612
rect 8412 19558 8458 19610
rect 8458 19558 8468 19610
rect 8492 19558 8522 19610
rect 8522 19558 8534 19610
rect 8534 19558 8548 19610
rect 8572 19558 8586 19610
rect 8586 19558 8598 19610
rect 8598 19558 8628 19610
rect 8652 19558 8662 19610
rect 8662 19558 8708 19610
rect 8412 19556 8468 19558
rect 8492 19556 8548 19558
rect 8572 19556 8628 19558
rect 8652 19556 8708 19558
rect 7752 19066 7808 19068
rect 7832 19066 7888 19068
rect 7912 19066 7968 19068
rect 7992 19066 8048 19068
rect 7752 19014 7798 19066
rect 7798 19014 7808 19066
rect 7832 19014 7862 19066
rect 7862 19014 7874 19066
rect 7874 19014 7888 19066
rect 7912 19014 7926 19066
rect 7926 19014 7938 19066
rect 7938 19014 7968 19066
rect 7992 19014 8002 19066
rect 8002 19014 8048 19066
rect 7752 19012 7808 19014
rect 7832 19012 7888 19014
rect 7912 19012 7968 19014
rect 7992 19012 8048 19014
rect 8412 18522 8468 18524
rect 8492 18522 8548 18524
rect 8572 18522 8628 18524
rect 8652 18522 8708 18524
rect 8412 18470 8458 18522
rect 8458 18470 8468 18522
rect 8492 18470 8522 18522
rect 8522 18470 8534 18522
rect 8534 18470 8548 18522
rect 8572 18470 8586 18522
rect 8586 18470 8598 18522
rect 8598 18470 8628 18522
rect 8652 18470 8662 18522
rect 8662 18470 8708 18522
rect 8412 18468 8468 18470
rect 8492 18468 8548 18470
rect 8572 18468 8628 18470
rect 8652 18468 8708 18470
rect 7752 17978 7808 17980
rect 7832 17978 7888 17980
rect 7912 17978 7968 17980
rect 7992 17978 8048 17980
rect 7752 17926 7798 17978
rect 7798 17926 7808 17978
rect 7832 17926 7862 17978
rect 7862 17926 7874 17978
rect 7874 17926 7888 17978
rect 7912 17926 7926 17978
rect 7926 17926 7938 17978
rect 7938 17926 7968 17978
rect 7992 17926 8002 17978
rect 8002 17926 8048 17978
rect 7752 17924 7808 17926
rect 7832 17924 7888 17926
rect 7912 17924 7968 17926
rect 7992 17924 8048 17926
rect 8412 17434 8468 17436
rect 8492 17434 8548 17436
rect 8572 17434 8628 17436
rect 8652 17434 8708 17436
rect 8412 17382 8458 17434
rect 8458 17382 8468 17434
rect 8492 17382 8522 17434
rect 8522 17382 8534 17434
rect 8534 17382 8548 17434
rect 8572 17382 8586 17434
rect 8586 17382 8598 17434
rect 8598 17382 8628 17434
rect 8652 17382 8662 17434
rect 8662 17382 8708 17434
rect 8412 17380 8468 17382
rect 8492 17380 8548 17382
rect 8572 17380 8628 17382
rect 8652 17380 8708 17382
rect 7752 16890 7808 16892
rect 7832 16890 7888 16892
rect 7912 16890 7968 16892
rect 7992 16890 8048 16892
rect 7752 16838 7798 16890
rect 7798 16838 7808 16890
rect 7832 16838 7862 16890
rect 7862 16838 7874 16890
rect 7874 16838 7888 16890
rect 7912 16838 7926 16890
rect 7926 16838 7938 16890
rect 7938 16838 7968 16890
rect 7992 16838 8002 16890
rect 8002 16838 8048 16890
rect 7752 16836 7808 16838
rect 7832 16836 7888 16838
rect 7912 16836 7968 16838
rect 7992 16836 8048 16838
rect 5262 12416 5318 12472
rect 5262 12280 5318 12336
rect 7752 15802 7808 15804
rect 7832 15802 7888 15804
rect 7912 15802 7968 15804
rect 7992 15802 8048 15804
rect 7752 15750 7798 15802
rect 7798 15750 7808 15802
rect 7832 15750 7862 15802
rect 7862 15750 7874 15802
rect 7874 15750 7888 15802
rect 7912 15750 7926 15802
rect 7926 15750 7938 15802
rect 7938 15750 7968 15802
rect 7992 15750 8002 15802
rect 8002 15750 8048 15802
rect 7752 15748 7808 15750
rect 7832 15748 7888 15750
rect 7912 15748 7968 15750
rect 7992 15748 8048 15750
rect 8412 16346 8468 16348
rect 8492 16346 8548 16348
rect 8572 16346 8628 16348
rect 8652 16346 8708 16348
rect 8412 16294 8458 16346
rect 8458 16294 8468 16346
rect 8492 16294 8522 16346
rect 8522 16294 8534 16346
rect 8534 16294 8548 16346
rect 8572 16294 8586 16346
rect 8586 16294 8598 16346
rect 8598 16294 8628 16346
rect 8652 16294 8662 16346
rect 8662 16294 8708 16346
rect 8412 16292 8468 16294
rect 8492 16292 8548 16294
rect 8572 16292 8628 16294
rect 8652 16292 8708 16294
rect 8412 15258 8468 15260
rect 8492 15258 8548 15260
rect 8572 15258 8628 15260
rect 8652 15258 8708 15260
rect 8412 15206 8458 15258
rect 8458 15206 8468 15258
rect 8492 15206 8522 15258
rect 8522 15206 8534 15258
rect 8534 15206 8548 15258
rect 8572 15206 8586 15258
rect 8586 15206 8598 15258
rect 8598 15206 8628 15258
rect 8652 15206 8662 15258
rect 8662 15206 8708 15258
rect 8412 15204 8468 15206
rect 8492 15204 8548 15206
rect 8572 15204 8628 15206
rect 8652 15204 8708 15206
rect 7752 14714 7808 14716
rect 7832 14714 7888 14716
rect 7912 14714 7968 14716
rect 7992 14714 8048 14716
rect 7752 14662 7798 14714
rect 7798 14662 7808 14714
rect 7832 14662 7862 14714
rect 7862 14662 7874 14714
rect 7874 14662 7888 14714
rect 7912 14662 7926 14714
rect 7926 14662 7938 14714
rect 7938 14662 7968 14714
rect 7992 14662 8002 14714
rect 8002 14662 8048 14714
rect 7752 14660 7808 14662
rect 7832 14660 7888 14662
rect 7912 14660 7968 14662
rect 7992 14660 8048 14662
rect 8412 14170 8468 14172
rect 8492 14170 8548 14172
rect 8572 14170 8628 14172
rect 8652 14170 8708 14172
rect 8412 14118 8458 14170
rect 8458 14118 8468 14170
rect 8492 14118 8522 14170
rect 8522 14118 8534 14170
rect 8534 14118 8548 14170
rect 8572 14118 8586 14170
rect 8586 14118 8598 14170
rect 8598 14118 8628 14170
rect 8652 14118 8662 14170
rect 8662 14118 8708 14170
rect 8412 14116 8468 14118
rect 8492 14116 8548 14118
rect 8572 14116 8628 14118
rect 8652 14116 8708 14118
rect 7752 13626 7808 13628
rect 7832 13626 7888 13628
rect 7912 13626 7968 13628
rect 7992 13626 8048 13628
rect 7752 13574 7798 13626
rect 7798 13574 7808 13626
rect 7832 13574 7862 13626
rect 7862 13574 7874 13626
rect 7874 13574 7888 13626
rect 7912 13574 7926 13626
rect 7926 13574 7938 13626
rect 7938 13574 7968 13626
rect 7992 13574 8002 13626
rect 8002 13574 8048 13626
rect 7752 13572 7808 13574
rect 7832 13572 7888 13574
rect 7912 13572 7968 13574
rect 7992 13572 8048 13574
rect 12283 20154 12339 20156
rect 12363 20154 12419 20156
rect 12443 20154 12499 20156
rect 12523 20154 12579 20156
rect 12283 20102 12329 20154
rect 12329 20102 12339 20154
rect 12363 20102 12393 20154
rect 12393 20102 12405 20154
rect 12405 20102 12419 20154
rect 12443 20102 12457 20154
rect 12457 20102 12469 20154
rect 12469 20102 12499 20154
rect 12523 20102 12533 20154
rect 12533 20102 12579 20154
rect 12283 20100 12339 20102
rect 12363 20100 12419 20102
rect 12443 20100 12499 20102
rect 12523 20100 12579 20102
rect 8412 13082 8468 13084
rect 8492 13082 8548 13084
rect 8572 13082 8628 13084
rect 8652 13082 8708 13084
rect 8412 13030 8458 13082
rect 8458 13030 8468 13082
rect 8492 13030 8522 13082
rect 8522 13030 8534 13082
rect 8534 13030 8548 13082
rect 8572 13030 8586 13082
rect 8586 13030 8598 13082
rect 8598 13030 8628 13082
rect 8652 13030 8662 13082
rect 8662 13030 8708 13082
rect 8412 13028 8468 13030
rect 8492 13028 8548 13030
rect 8572 13028 8628 13030
rect 8652 13028 8708 13030
rect 7752 12538 7808 12540
rect 7832 12538 7888 12540
rect 7912 12538 7968 12540
rect 7992 12538 8048 12540
rect 7752 12486 7798 12538
rect 7798 12486 7808 12538
rect 7832 12486 7862 12538
rect 7862 12486 7874 12538
rect 7874 12486 7888 12538
rect 7912 12486 7926 12538
rect 7926 12486 7938 12538
rect 7938 12486 7968 12538
rect 7992 12486 8002 12538
rect 8002 12486 8048 12538
rect 7752 12484 7808 12486
rect 7832 12484 7888 12486
rect 7912 12484 7968 12486
rect 7992 12484 8048 12486
rect 8412 11994 8468 11996
rect 8492 11994 8548 11996
rect 8572 11994 8628 11996
rect 8652 11994 8708 11996
rect 8412 11942 8458 11994
rect 8458 11942 8468 11994
rect 8492 11942 8522 11994
rect 8522 11942 8534 11994
rect 8534 11942 8548 11994
rect 8572 11942 8586 11994
rect 8586 11942 8598 11994
rect 8598 11942 8628 11994
rect 8652 11942 8662 11994
rect 8662 11942 8708 11994
rect 8412 11940 8468 11942
rect 8492 11940 8548 11942
rect 8572 11940 8628 11942
rect 8652 11940 8708 11942
rect 7752 11450 7808 11452
rect 7832 11450 7888 11452
rect 7912 11450 7968 11452
rect 7992 11450 8048 11452
rect 7752 11398 7798 11450
rect 7798 11398 7808 11450
rect 7832 11398 7862 11450
rect 7862 11398 7874 11450
rect 7874 11398 7888 11450
rect 7912 11398 7926 11450
rect 7926 11398 7938 11450
rect 7938 11398 7968 11450
rect 7992 11398 8002 11450
rect 8002 11398 8048 11450
rect 7752 11396 7808 11398
rect 7832 11396 7888 11398
rect 7912 11396 7968 11398
rect 7992 11396 8048 11398
rect 8412 10906 8468 10908
rect 8492 10906 8548 10908
rect 8572 10906 8628 10908
rect 8652 10906 8708 10908
rect 8412 10854 8458 10906
rect 8458 10854 8468 10906
rect 8492 10854 8522 10906
rect 8522 10854 8534 10906
rect 8534 10854 8548 10906
rect 8572 10854 8586 10906
rect 8586 10854 8598 10906
rect 8598 10854 8628 10906
rect 8652 10854 8662 10906
rect 8662 10854 8708 10906
rect 8412 10852 8468 10854
rect 8492 10852 8548 10854
rect 8572 10852 8628 10854
rect 8652 10852 8708 10854
rect 7752 10362 7808 10364
rect 7832 10362 7888 10364
rect 7912 10362 7968 10364
rect 7992 10362 8048 10364
rect 7752 10310 7798 10362
rect 7798 10310 7808 10362
rect 7832 10310 7862 10362
rect 7862 10310 7874 10362
rect 7874 10310 7888 10362
rect 7912 10310 7926 10362
rect 7926 10310 7938 10362
rect 7938 10310 7968 10362
rect 7992 10310 8002 10362
rect 8002 10310 8048 10362
rect 7752 10308 7808 10310
rect 7832 10308 7888 10310
rect 7912 10308 7968 10310
rect 7992 10308 8048 10310
rect 9770 12300 9826 12336
rect 9770 12280 9772 12300
rect 9772 12280 9824 12300
rect 9824 12280 9826 12300
rect 8412 9818 8468 9820
rect 8492 9818 8548 9820
rect 8572 9818 8628 9820
rect 8652 9818 8708 9820
rect 8412 9766 8458 9818
rect 8458 9766 8468 9818
rect 8492 9766 8522 9818
rect 8522 9766 8534 9818
rect 8534 9766 8548 9818
rect 8572 9766 8586 9818
rect 8586 9766 8598 9818
rect 8598 9766 8628 9818
rect 8652 9766 8662 9818
rect 8662 9766 8708 9818
rect 8412 9764 8468 9766
rect 8492 9764 8548 9766
rect 8572 9764 8628 9766
rect 8652 9764 8708 9766
rect 7752 9274 7808 9276
rect 7832 9274 7888 9276
rect 7912 9274 7968 9276
rect 7992 9274 8048 9276
rect 7752 9222 7798 9274
rect 7798 9222 7808 9274
rect 7832 9222 7862 9274
rect 7862 9222 7874 9274
rect 7874 9222 7888 9274
rect 7912 9222 7926 9274
rect 7926 9222 7938 9274
rect 7938 9222 7968 9274
rect 7992 9222 8002 9274
rect 8002 9222 8048 9274
rect 7752 9220 7808 9222
rect 7832 9220 7888 9222
rect 7912 9220 7968 9222
rect 7992 9220 8048 9222
rect 3221 7098 3277 7100
rect 3301 7098 3357 7100
rect 3381 7098 3437 7100
rect 3461 7098 3517 7100
rect 3221 7046 3267 7098
rect 3267 7046 3277 7098
rect 3301 7046 3331 7098
rect 3331 7046 3343 7098
rect 3343 7046 3357 7098
rect 3381 7046 3395 7098
rect 3395 7046 3407 7098
rect 3407 7046 3437 7098
rect 3461 7046 3471 7098
rect 3471 7046 3517 7098
rect 3221 7044 3277 7046
rect 3301 7044 3357 7046
rect 3381 7044 3437 7046
rect 3461 7044 3517 7046
rect 3881 6554 3937 6556
rect 3961 6554 4017 6556
rect 4041 6554 4097 6556
rect 4121 6554 4177 6556
rect 3881 6502 3927 6554
rect 3927 6502 3937 6554
rect 3961 6502 3991 6554
rect 3991 6502 4003 6554
rect 4003 6502 4017 6554
rect 4041 6502 4055 6554
rect 4055 6502 4067 6554
rect 4067 6502 4097 6554
rect 4121 6502 4131 6554
rect 4131 6502 4177 6554
rect 3881 6500 3937 6502
rect 3961 6500 4017 6502
rect 4041 6500 4097 6502
rect 4121 6500 4177 6502
rect 3221 6010 3277 6012
rect 3301 6010 3357 6012
rect 3381 6010 3437 6012
rect 3461 6010 3517 6012
rect 3221 5958 3267 6010
rect 3267 5958 3277 6010
rect 3301 5958 3331 6010
rect 3331 5958 3343 6010
rect 3343 5958 3357 6010
rect 3381 5958 3395 6010
rect 3395 5958 3407 6010
rect 3407 5958 3437 6010
rect 3461 5958 3471 6010
rect 3471 5958 3517 6010
rect 3221 5956 3277 5958
rect 3301 5956 3357 5958
rect 3381 5956 3437 5958
rect 3461 5956 3517 5958
rect 8412 8730 8468 8732
rect 8492 8730 8548 8732
rect 8572 8730 8628 8732
rect 8652 8730 8708 8732
rect 8412 8678 8458 8730
rect 8458 8678 8468 8730
rect 8492 8678 8522 8730
rect 8522 8678 8534 8730
rect 8534 8678 8548 8730
rect 8572 8678 8586 8730
rect 8586 8678 8598 8730
rect 8598 8678 8628 8730
rect 8652 8678 8662 8730
rect 8662 8678 8708 8730
rect 8412 8676 8468 8678
rect 8492 8676 8548 8678
rect 8572 8676 8628 8678
rect 8652 8676 8708 8678
rect 7752 8186 7808 8188
rect 7832 8186 7888 8188
rect 7912 8186 7968 8188
rect 7992 8186 8048 8188
rect 7752 8134 7798 8186
rect 7798 8134 7808 8186
rect 7832 8134 7862 8186
rect 7862 8134 7874 8186
rect 7874 8134 7888 8186
rect 7912 8134 7926 8186
rect 7926 8134 7938 8186
rect 7938 8134 7968 8186
rect 7992 8134 8002 8186
rect 8002 8134 8048 8186
rect 7752 8132 7808 8134
rect 7832 8132 7888 8134
rect 7912 8132 7968 8134
rect 7992 8132 8048 8134
rect 3221 4922 3277 4924
rect 3301 4922 3357 4924
rect 3381 4922 3437 4924
rect 3461 4922 3517 4924
rect 3221 4870 3267 4922
rect 3267 4870 3277 4922
rect 3301 4870 3331 4922
rect 3331 4870 3343 4922
rect 3343 4870 3357 4922
rect 3381 4870 3395 4922
rect 3395 4870 3407 4922
rect 3407 4870 3437 4922
rect 3461 4870 3471 4922
rect 3471 4870 3517 4922
rect 3221 4868 3277 4870
rect 3301 4868 3357 4870
rect 3381 4868 3437 4870
rect 3461 4868 3517 4870
rect 3881 5466 3937 5468
rect 3961 5466 4017 5468
rect 4041 5466 4097 5468
rect 4121 5466 4177 5468
rect 3881 5414 3927 5466
rect 3927 5414 3937 5466
rect 3961 5414 3991 5466
rect 3991 5414 4003 5466
rect 4003 5414 4017 5466
rect 4041 5414 4055 5466
rect 4055 5414 4067 5466
rect 4067 5414 4097 5466
rect 4121 5414 4131 5466
rect 4131 5414 4177 5466
rect 3881 5412 3937 5414
rect 3961 5412 4017 5414
rect 4041 5412 4097 5414
rect 4121 5412 4177 5414
rect 8412 7642 8468 7644
rect 8492 7642 8548 7644
rect 8572 7642 8628 7644
rect 8652 7642 8708 7644
rect 8412 7590 8458 7642
rect 8458 7590 8468 7642
rect 8492 7590 8522 7642
rect 8522 7590 8534 7642
rect 8534 7590 8548 7642
rect 8572 7590 8586 7642
rect 8586 7590 8598 7642
rect 8598 7590 8628 7642
rect 8652 7590 8662 7642
rect 8662 7590 8708 7642
rect 8412 7588 8468 7590
rect 8492 7588 8548 7590
rect 8572 7588 8628 7590
rect 8652 7588 8708 7590
rect 7752 7098 7808 7100
rect 7832 7098 7888 7100
rect 7912 7098 7968 7100
rect 7992 7098 8048 7100
rect 7752 7046 7798 7098
rect 7798 7046 7808 7098
rect 7832 7046 7862 7098
rect 7862 7046 7874 7098
rect 7874 7046 7888 7098
rect 7912 7046 7926 7098
rect 7926 7046 7938 7098
rect 7938 7046 7968 7098
rect 7992 7046 8002 7098
rect 8002 7046 8048 7098
rect 7752 7044 7808 7046
rect 7832 7044 7888 7046
rect 7912 7044 7968 7046
rect 7992 7044 8048 7046
rect 8412 6554 8468 6556
rect 8492 6554 8548 6556
rect 8572 6554 8628 6556
rect 8652 6554 8708 6556
rect 8412 6502 8458 6554
rect 8458 6502 8468 6554
rect 8492 6502 8522 6554
rect 8522 6502 8534 6554
rect 8534 6502 8548 6554
rect 8572 6502 8586 6554
rect 8586 6502 8598 6554
rect 8598 6502 8628 6554
rect 8652 6502 8662 6554
rect 8662 6502 8708 6554
rect 8412 6500 8468 6502
rect 8492 6500 8548 6502
rect 8572 6500 8628 6502
rect 8652 6500 8708 6502
rect 7752 6010 7808 6012
rect 7832 6010 7888 6012
rect 7912 6010 7968 6012
rect 7992 6010 8048 6012
rect 7752 5958 7798 6010
rect 7798 5958 7808 6010
rect 7832 5958 7862 6010
rect 7862 5958 7874 6010
rect 7874 5958 7888 6010
rect 7912 5958 7926 6010
rect 7926 5958 7938 6010
rect 7938 5958 7968 6010
rect 7992 5958 8002 6010
rect 8002 5958 8048 6010
rect 7752 5956 7808 5958
rect 7832 5956 7888 5958
rect 7912 5956 7968 5958
rect 7992 5956 8048 5958
rect 11058 11192 11114 11248
rect 12943 19610 12999 19612
rect 13023 19610 13079 19612
rect 13103 19610 13159 19612
rect 13183 19610 13239 19612
rect 12943 19558 12989 19610
rect 12989 19558 12999 19610
rect 13023 19558 13053 19610
rect 13053 19558 13065 19610
rect 13065 19558 13079 19610
rect 13103 19558 13117 19610
rect 13117 19558 13129 19610
rect 13129 19558 13159 19610
rect 13183 19558 13193 19610
rect 13193 19558 13239 19610
rect 12943 19556 12999 19558
rect 13023 19556 13079 19558
rect 13103 19556 13159 19558
rect 13183 19556 13239 19558
rect 12283 19066 12339 19068
rect 12363 19066 12419 19068
rect 12443 19066 12499 19068
rect 12523 19066 12579 19068
rect 12283 19014 12329 19066
rect 12329 19014 12339 19066
rect 12363 19014 12393 19066
rect 12393 19014 12405 19066
rect 12405 19014 12419 19066
rect 12443 19014 12457 19066
rect 12457 19014 12469 19066
rect 12469 19014 12499 19066
rect 12523 19014 12533 19066
rect 12533 19014 12579 19066
rect 12283 19012 12339 19014
rect 12363 19012 12419 19014
rect 12443 19012 12499 19014
rect 12523 19012 12579 19014
rect 12943 18522 12999 18524
rect 13023 18522 13079 18524
rect 13103 18522 13159 18524
rect 13183 18522 13239 18524
rect 12943 18470 12989 18522
rect 12989 18470 12999 18522
rect 13023 18470 13053 18522
rect 13053 18470 13065 18522
rect 13065 18470 13079 18522
rect 13103 18470 13117 18522
rect 13117 18470 13129 18522
rect 13129 18470 13159 18522
rect 13183 18470 13193 18522
rect 13193 18470 13239 18522
rect 12943 18468 12999 18470
rect 13023 18468 13079 18470
rect 13103 18468 13159 18470
rect 13183 18468 13239 18470
rect 12283 17978 12339 17980
rect 12363 17978 12419 17980
rect 12443 17978 12499 17980
rect 12523 17978 12579 17980
rect 12283 17926 12329 17978
rect 12329 17926 12339 17978
rect 12363 17926 12393 17978
rect 12393 17926 12405 17978
rect 12405 17926 12419 17978
rect 12443 17926 12457 17978
rect 12457 17926 12469 17978
rect 12469 17926 12499 17978
rect 12523 17926 12533 17978
rect 12533 17926 12579 17978
rect 12283 17924 12339 17926
rect 12363 17924 12419 17926
rect 12443 17924 12499 17926
rect 12523 17924 12579 17926
rect 12943 17434 12999 17436
rect 13023 17434 13079 17436
rect 13103 17434 13159 17436
rect 13183 17434 13239 17436
rect 12943 17382 12989 17434
rect 12989 17382 12999 17434
rect 13023 17382 13053 17434
rect 13053 17382 13065 17434
rect 13065 17382 13079 17434
rect 13103 17382 13117 17434
rect 13117 17382 13129 17434
rect 13129 17382 13159 17434
rect 13183 17382 13193 17434
rect 13193 17382 13239 17434
rect 12943 17380 12999 17382
rect 13023 17380 13079 17382
rect 13103 17380 13159 17382
rect 13183 17380 13239 17382
rect 12283 16890 12339 16892
rect 12363 16890 12419 16892
rect 12443 16890 12499 16892
rect 12523 16890 12579 16892
rect 12283 16838 12329 16890
rect 12329 16838 12339 16890
rect 12363 16838 12393 16890
rect 12393 16838 12405 16890
rect 12405 16838 12419 16890
rect 12443 16838 12457 16890
rect 12457 16838 12469 16890
rect 12469 16838 12499 16890
rect 12523 16838 12533 16890
rect 12533 16838 12579 16890
rect 12283 16836 12339 16838
rect 12363 16836 12419 16838
rect 12443 16836 12499 16838
rect 12523 16836 12579 16838
rect 12943 16346 12999 16348
rect 13023 16346 13079 16348
rect 13103 16346 13159 16348
rect 13183 16346 13239 16348
rect 12943 16294 12989 16346
rect 12989 16294 12999 16346
rect 13023 16294 13053 16346
rect 13053 16294 13065 16346
rect 13065 16294 13079 16346
rect 13103 16294 13117 16346
rect 13117 16294 13129 16346
rect 13129 16294 13159 16346
rect 13183 16294 13193 16346
rect 13193 16294 13239 16346
rect 12943 16292 12999 16294
rect 13023 16292 13079 16294
rect 13103 16292 13159 16294
rect 13183 16292 13239 16294
rect 12283 15802 12339 15804
rect 12363 15802 12419 15804
rect 12443 15802 12499 15804
rect 12523 15802 12579 15804
rect 12283 15750 12329 15802
rect 12329 15750 12339 15802
rect 12363 15750 12393 15802
rect 12393 15750 12405 15802
rect 12405 15750 12419 15802
rect 12443 15750 12457 15802
rect 12457 15750 12469 15802
rect 12469 15750 12499 15802
rect 12523 15750 12533 15802
rect 12533 15750 12579 15802
rect 12283 15748 12339 15750
rect 12363 15748 12419 15750
rect 12443 15748 12499 15750
rect 12523 15748 12579 15750
rect 12943 15258 12999 15260
rect 13023 15258 13079 15260
rect 13103 15258 13159 15260
rect 13183 15258 13239 15260
rect 12943 15206 12989 15258
rect 12989 15206 12999 15258
rect 13023 15206 13053 15258
rect 13053 15206 13065 15258
rect 13065 15206 13079 15258
rect 13103 15206 13117 15258
rect 13117 15206 13129 15258
rect 13129 15206 13159 15258
rect 13183 15206 13193 15258
rect 13193 15206 13239 15258
rect 12943 15204 12999 15206
rect 13023 15204 13079 15206
rect 13103 15204 13159 15206
rect 13183 15204 13239 15206
rect 12283 14714 12339 14716
rect 12363 14714 12419 14716
rect 12443 14714 12499 14716
rect 12523 14714 12579 14716
rect 12283 14662 12329 14714
rect 12329 14662 12339 14714
rect 12363 14662 12393 14714
rect 12393 14662 12405 14714
rect 12405 14662 12419 14714
rect 12443 14662 12457 14714
rect 12457 14662 12469 14714
rect 12469 14662 12499 14714
rect 12523 14662 12533 14714
rect 12533 14662 12579 14714
rect 12283 14660 12339 14662
rect 12363 14660 12419 14662
rect 12443 14660 12499 14662
rect 12523 14660 12579 14662
rect 12943 14170 12999 14172
rect 13023 14170 13079 14172
rect 13103 14170 13159 14172
rect 13183 14170 13239 14172
rect 12943 14118 12989 14170
rect 12989 14118 12999 14170
rect 13023 14118 13053 14170
rect 13053 14118 13065 14170
rect 13065 14118 13079 14170
rect 13103 14118 13117 14170
rect 13117 14118 13129 14170
rect 13129 14118 13159 14170
rect 13183 14118 13193 14170
rect 13193 14118 13239 14170
rect 12943 14116 12999 14118
rect 13023 14116 13079 14118
rect 13103 14116 13159 14118
rect 13183 14116 13239 14118
rect 12283 13626 12339 13628
rect 12363 13626 12419 13628
rect 12443 13626 12499 13628
rect 12523 13626 12579 13628
rect 12283 13574 12329 13626
rect 12329 13574 12339 13626
rect 12363 13574 12393 13626
rect 12393 13574 12405 13626
rect 12405 13574 12419 13626
rect 12443 13574 12457 13626
rect 12457 13574 12469 13626
rect 12469 13574 12499 13626
rect 12523 13574 12533 13626
rect 12533 13574 12579 13626
rect 12283 13572 12339 13574
rect 12363 13572 12419 13574
rect 12443 13572 12499 13574
rect 12523 13572 12579 13574
rect 12943 13082 12999 13084
rect 13023 13082 13079 13084
rect 13103 13082 13159 13084
rect 13183 13082 13239 13084
rect 12943 13030 12989 13082
rect 12989 13030 12999 13082
rect 13023 13030 13053 13082
rect 13053 13030 13065 13082
rect 13065 13030 13079 13082
rect 13103 13030 13117 13082
rect 13117 13030 13129 13082
rect 13129 13030 13159 13082
rect 13183 13030 13193 13082
rect 13193 13030 13239 13082
rect 12943 13028 12999 13030
rect 13023 13028 13079 13030
rect 13103 13028 13159 13030
rect 13183 13028 13239 13030
rect 12283 12538 12339 12540
rect 12363 12538 12419 12540
rect 12443 12538 12499 12540
rect 12523 12538 12579 12540
rect 12283 12486 12329 12538
rect 12329 12486 12339 12538
rect 12363 12486 12393 12538
rect 12393 12486 12405 12538
rect 12405 12486 12419 12538
rect 12443 12486 12457 12538
rect 12457 12486 12469 12538
rect 12469 12486 12499 12538
rect 12523 12486 12533 12538
rect 12533 12486 12579 12538
rect 12283 12484 12339 12486
rect 12363 12484 12419 12486
rect 12443 12484 12499 12486
rect 12523 12484 12579 12486
rect 12806 12280 12862 12336
rect 12283 11450 12339 11452
rect 12363 11450 12419 11452
rect 12443 11450 12499 11452
rect 12523 11450 12579 11452
rect 12283 11398 12329 11450
rect 12329 11398 12339 11450
rect 12363 11398 12393 11450
rect 12393 11398 12405 11450
rect 12405 11398 12419 11450
rect 12443 11398 12457 11450
rect 12457 11398 12469 11450
rect 12469 11398 12499 11450
rect 12523 11398 12533 11450
rect 12533 11398 12579 11450
rect 12283 11396 12339 11398
rect 12363 11396 12419 11398
rect 12443 11396 12499 11398
rect 12523 11396 12579 11398
rect 12283 10362 12339 10364
rect 12363 10362 12419 10364
rect 12443 10362 12499 10364
rect 12523 10362 12579 10364
rect 12283 10310 12329 10362
rect 12329 10310 12339 10362
rect 12363 10310 12393 10362
rect 12393 10310 12405 10362
rect 12405 10310 12419 10362
rect 12443 10310 12457 10362
rect 12457 10310 12469 10362
rect 12469 10310 12499 10362
rect 12523 10310 12533 10362
rect 12533 10310 12579 10362
rect 12283 10308 12339 10310
rect 12363 10308 12419 10310
rect 12443 10308 12499 10310
rect 12523 10308 12579 10310
rect 12283 9274 12339 9276
rect 12363 9274 12419 9276
rect 12443 9274 12499 9276
rect 12523 9274 12579 9276
rect 12283 9222 12329 9274
rect 12329 9222 12339 9274
rect 12363 9222 12393 9274
rect 12393 9222 12405 9274
rect 12405 9222 12419 9274
rect 12443 9222 12457 9274
rect 12457 9222 12469 9274
rect 12469 9222 12499 9274
rect 12523 9222 12533 9274
rect 12533 9222 12579 9274
rect 12283 9220 12339 9222
rect 12363 9220 12419 9222
rect 12443 9220 12499 9222
rect 12523 9220 12579 9222
rect 12943 11994 12999 11996
rect 13023 11994 13079 11996
rect 13103 11994 13159 11996
rect 13183 11994 13239 11996
rect 12943 11942 12989 11994
rect 12989 11942 12999 11994
rect 13023 11942 13053 11994
rect 13053 11942 13065 11994
rect 13065 11942 13079 11994
rect 13103 11942 13117 11994
rect 13117 11942 13129 11994
rect 13129 11942 13159 11994
rect 13183 11942 13193 11994
rect 13193 11942 13239 11994
rect 12943 11940 12999 11942
rect 13023 11940 13079 11942
rect 13103 11940 13159 11942
rect 13183 11940 13239 11942
rect 12943 10906 12999 10908
rect 13023 10906 13079 10908
rect 13103 10906 13159 10908
rect 13183 10906 13239 10908
rect 12943 10854 12989 10906
rect 12989 10854 12999 10906
rect 13023 10854 13053 10906
rect 13053 10854 13065 10906
rect 13065 10854 13079 10906
rect 13103 10854 13117 10906
rect 13117 10854 13129 10906
rect 13129 10854 13159 10906
rect 13183 10854 13193 10906
rect 13193 10854 13239 10906
rect 12943 10852 12999 10854
rect 13023 10852 13079 10854
rect 13103 10852 13159 10854
rect 13183 10852 13239 10854
rect 12943 9818 12999 9820
rect 13023 9818 13079 9820
rect 13103 9818 13159 9820
rect 13183 9818 13239 9820
rect 12943 9766 12989 9818
rect 12989 9766 12999 9818
rect 13023 9766 13053 9818
rect 13053 9766 13065 9818
rect 13065 9766 13079 9818
rect 13103 9766 13117 9818
rect 13117 9766 13129 9818
rect 13129 9766 13159 9818
rect 13183 9766 13193 9818
rect 13193 9766 13239 9818
rect 12943 9764 12999 9766
rect 13023 9764 13079 9766
rect 13103 9764 13159 9766
rect 13183 9764 13239 9766
rect 16814 20154 16870 20156
rect 16894 20154 16950 20156
rect 16974 20154 17030 20156
rect 17054 20154 17110 20156
rect 16814 20102 16860 20154
rect 16860 20102 16870 20154
rect 16894 20102 16924 20154
rect 16924 20102 16936 20154
rect 16936 20102 16950 20154
rect 16974 20102 16988 20154
rect 16988 20102 17000 20154
rect 17000 20102 17030 20154
rect 17054 20102 17064 20154
rect 17064 20102 17110 20154
rect 16814 20100 16870 20102
rect 16894 20100 16950 20102
rect 16974 20100 17030 20102
rect 17054 20100 17110 20102
rect 12943 8730 12999 8732
rect 13023 8730 13079 8732
rect 13103 8730 13159 8732
rect 13183 8730 13239 8732
rect 12943 8678 12989 8730
rect 12989 8678 12999 8730
rect 13023 8678 13053 8730
rect 13053 8678 13065 8730
rect 13065 8678 13079 8730
rect 13103 8678 13117 8730
rect 13117 8678 13129 8730
rect 13129 8678 13159 8730
rect 13183 8678 13193 8730
rect 13193 8678 13239 8730
rect 12943 8676 12999 8678
rect 13023 8676 13079 8678
rect 13103 8676 13159 8678
rect 13183 8676 13239 8678
rect 12283 8186 12339 8188
rect 12363 8186 12419 8188
rect 12443 8186 12499 8188
rect 12523 8186 12579 8188
rect 12283 8134 12329 8186
rect 12329 8134 12339 8186
rect 12363 8134 12393 8186
rect 12393 8134 12405 8186
rect 12405 8134 12419 8186
rect 12443 8134 12457 8186
rect 12457 8134 12469 8186
rect 12469 8134 12499 8186
rect 12523 8134 12533 8186
rect 12533 8134 12579 8186
rect 12283 8132 12339 8134
rect 12363 8132 12419 8134
rect 12443 8132 12499 8134
rect 12523 8132 12579 8134
rect 8412 5466 8468 5468
rect 8492 5466 8548 5468
rect 8572 5466 8628 5468
rect 8652 5466 8708 5468
rect 8412 5414 8458 5466
rect 8458 5414 8468 5466
rect 8492 5414 8522 5466
rect 8522 5414 8534 5466
rect 8534 5414 8548 5466
rect 8572 5414 8586 5466
rect 8586 5414 8598 5466
rect 8598 5414 8628 5466
rect 8652 5414 8662 5466
rect 8662 5414 8708 5466
rect 8412 5412 8468 5414
rect 8492 5412 8548 5414
rect 8572 5412 8628 5414
rect 8652 5412 8708 5414
rect 12943 7642 12999 7644
rect 13023 7642 13079 7644
rect 13103 7642 13159 7644
rect 13183 7642 13239 7644
rect 12943 7590 12989 7642
rect 12989 7590 12999 7642
rect 13023 7590 13053 7642
rect 13053 7590 13065 7642
rect 13065 7590 13079 7642
rect 13103 7590 13117 7642
rect 13117 7590 13129 7642
rect 13129 7590 13159 7642
rect 13183 7590 13193 7642
rect 13193 7590 13239 7642
rect 12943 7588 12999 7590
rect 13023 7588 13079 7590
rect 13103 7588 13159 7590
rect 13183 7588 13239 7590
rect 12283 7098 12339 7100
rect 12363 7098 12419 7100
rect 12443 7098 12499 7100
rect 12523 7098 12579 7100
rect 12283 7046 12329 7098
rect 12329 7046 12339 7098
rect 12363 7046 12393 7098
rect 12393 7046 12405 7098
rect 12405 7046 12419 7098
rect 12443 7046 12457 7098
rect 12457 7046 12469 7098
rect 12469 7046 12499 7098
rect 12523 7046 12533 7098
rect 12533 7046 12579 7098
rect 12283 7044 12339 7046
rect 12363 7044 12419 7046
rect 12443 7044 12499 7046
rect 12523 7044 12579 7046
rect 12283 6010 12339 6012
rect 12363 6010 12419 6012
rect 12443 6010 12499 6012
rect 12523 6010 12579 6012
rect 12283 5958 12329 6010
rect 12329 5958 12339 6010
rect 12363 5958 12393 6010
rect 12393 5958 12405 6010
rect 12405 5958 12419 6010
rect 12443 5958 12457 6010
rect 12457 5958 12469 6010
rect 12469 5958 12499 6010
rect 12523 5958 12533 6010
rect 12533 5958 12579 6010
rect 12283 5956 12339 5958
rect 12363 5956 12419 5958
rect 12443 5956 12499 5958
rect 12523 5956 12579 5958
rect 7752 4922 7808 4924
rect 7832 4922 7888 4924
rect 7912 4922 7968 4924
rect 7992 4922 8048 4924
rect 7752 4870 7798 4922
rect 7798 4870 7808 4922
rect 7832 4870 7862 4922
rect 7862 4870 7874 4922
rect 7874 4870 7888 4922
rect 7912 4870 7926 4922
rect 7926 4870 7938 4922
rect 7938 4870 7968 4922
rect 7992 4870 8002 4922
rect 8002 4870 8048 4922
rect 7752 4868 7808 4870
rect 7832 4868 7888 4870
rect 7912 4868 7968 4870
rect 7992 4868 8048 4870
rect 12943 6554 12999 6556
rect 13023 6554 13079 6556
rect 13103 6554 13159 6556
rect 13183 6554 13239 6556
rect 12943 6502 12989 6554
rect 12989 6502 12999 6554
rect 13023 6502 13053 6554
rect 13053 6502 13065 6554
rect 13065 6502 13079 6554
rect 13103 6502 13117 6554
rect 13117 6502 13129 6554
rect 13129 6502 13159 6554
rect 13183 6502 13193 6554
rect 13193 6502 13239 6554
rect 12943 6500 12999 6502
rect 13023 6500 13079 6502
rect 13103 6500 13159 6502
rect 13183 6500 13239 6502
rect 12283 4922 12339 4924
rect 12363 4922 12419 4924
rect 12443 4922 12499 4924
rect 12523 4922 12579 4924
rect 12283 4870 12329 4922
rect 12329 4870 12339 4922
rect 12363 4870 12393 4922
rect 12393 4870 12405 4922
rect 12405 4870 12419 4922
rect 12443 4870 12457 4922
rect 12457 4870 12469 4922
rect 12469 4870 12499 4922
rect 12523 4870 12533 4922
rect 12533 4870 12579 4922
rect 12283 4868 12339 4870
rect 12363 4868 12419 4870
rect 12443 4868 12499 4870
rect 12523 4868 12579 4870
rect 12943 5466 12999 5468
rect 13023 5466 13079 5468
rect 13103 5466 13159 5468
rect 13183 5466 13239 5468
rect 12943 5414 12989 5466
rect 12989 5414 12999 5466
rect 13023 5414 13053 5466
rect 13053 5414 13065 5466
rect 13065 5414 13079 5466
rect 13103 5414 13117 5466
rect 13117 5414 13129 5466
rect 13129 5414 13159 5466
rect 13183 5414 13193 5466
rect 13193 5414 13239 5466
rect 12943 5412 12999 5414
rect 13023 5412 13079 5414
rect 13103 5412 13159 5414
rect 13183 5412 13239 5414
rect 17130 19760 17186 19816
rect 16814 19066 16870 19068
rect 16894 19066 16950 19068
rect 16974 19066 17030 19068
rect 17054 19066 17110 19068
rect 16814 19014 16860 19066
rect 16860 19014 16870 19066
rect 16894 19014 16924 19066
rect 16924 19014 16936 19066
rect 16936 19014 16950 19066
rect 16974 19014 16988 19066
rect 16988 19014 17000 19066
rect 17000 19014 17030 19066
rect 17054 19014 17064 19066
rect 17064 19014 17110 19066
rect 16814 19012 16870 19014
rect 16894 19012 16950 19014
rect 16974 19012 17030 19014
rect 17054 19012 17110 19014
rect 16814 17978 16870 17980
rect 16894 17978 16950 17980
rect 16974 17978 17030 17980
rect 17054 17978 17110 17980
rect 16814 17926 16860 17978
rect 16860 17926 16870 17978
rect 16894 17926 16924 17978
rect 16924 17926 16936 17978
rect 16936 17926 16950 17978
rect 16974 17926 16988 17978
rect 16988 17926 17000 17978
rect 17000 17926 17030 17978
rect 17054 17926 17064 17978
rect 17064 17926 17110 17978
rect 16814 17924 16870 17926
rect 16894 17924 16950 17926
rect 16974 17924 17030 17926
rect 17054 17924 17110 17926
rect 16814 16890 16870 16892
rect 16894 16890 16950 16892
rect 16974 16890 17030 16892
rect 17054 16890 17110 16892
rect 16814 16838 16860 16890
rect 16860 16838 16870 16890
rect 16894 16838 16924 16890
rect 16924 16838 16936 16890
rect 16936 16838 16950 16890
rect 16974 16838 16988 16890
rect 16988 16838 17000 16890
rect 17000 16838 17030 16890
rect 17054 16838 17064 16890
rect 17064 16838 17110 16890
rect 16814 16836 16870 16838
rect 16894 16836 16950 16838
rect 16974 16836 17030 16838
rect 17054 16836 17110 16838
rect 16814 15802 16870 15804
rect 16894 15802 16950 15804
rect 16974 15802 17030 15804
rect 17054 15802 17110 15804
rect 16814 15750 16860 15802
rect 16860 15750 16870 15802
rect 16894 15750 16924 15802
rect 16924 15750 16936 15802
rect 16936 15750 16950 15802
rect 16974 15750 16988 15802
rect 16988 15750 17000 15802
rect 17000 15750 17030 15802
rect 17054 15750 17064 15802
rect 17064 15750 17110 15802
rect 16814 15748 16870 15750
rect 16894 15748 16950 15750
rect 16974 15748 17030 15750
rect 17054 15748 17110 15750
rect 16814 14714 16870 14716
rect 16894 14714 16950 14716
rect 16974 14714 17030 14716
rect 17054 14714 17110 14716
rect 16814 14662 16860 14714
rect 16860 14662 16870 14714
rect 16894 14662 16924 14714
rect 16924 14662 16936 14714
rect 16936 14662 16950 14714
rect 16974 14662 16988 14714
rect 16988 14662 17000 14714
rect 17000 14662 17030 14714
rect 17054 14662 17064 14714
rect 17064 14662 17110 14714
rect 16814 14660 16870 14662
rect 16894 14660 16950 14662
rect 16974 14660 17030 14662
rect 17054 14660 17110 14662
rect 17682 19760 17738 19816
rect 17474 19610 17530 19612
rect 17554 19610 17610 19612
rect 17634 19610 17690 19612
rect 17714 19610 17770 19612
rect 17474 19558 17520 19610
rect 17520 19558 17530 19610
rect 17554 19558 17584 19610
rect 17584 19558 17596 19610
rect 17596 19558 17610 19610
rect 17634 19558 17648 19610
rect 17648 19558 17660 19610
rect 17660 19558 17690 19610
rect 17714 19558 17724 19610
rect 17724 19558 17770 19610
rect 17474 19556 17530 19558
rect 17554 19556 17610 19558
rect 17634 19556 17690 19558
rect 17714 19556 17770 19558
rect 17474 18522 17530 18524
rect 17554 18522 17610 18524
rect 17634 18522 17690 18524
rect 17714 18522 17770 18524
rect 17474 18470 17520 18522
rect 17520 18470 17530 18522
rect 17554 18470 17584 18522
rect 17584 18470 17596 18522
rect 17596 18470 17610 18522
rect 17634 18470 17648 18522
rect 17648 18470 17660 18522
rect 17660 18470 17690 18522
rect 17714 18470 17724 18522
rect 17724 18470 17770 18522
rect 17474 18468 17530 18470
rect 17554 18468 17610 18470
rect 17634 18468 17690 18470
rect 17714 18468 17770 18470
rect 17474 17434 17530 17436
rect 17554 17434 17610 17436
rect 17634 17434 17690 17436
rect 17714 17434 17770 17436
rect 17474 17382 17520 17434
rect 17520 17382 17530 17434
rect 17554 17382 17584 17434
rect 17584 17382 17596 17434
rect 17596 17382 17610 17434
rect 17634 17382 17648 17434
rect 17648 17382 17660 17434
rect 17660 17382 17690 17434
rect 17714 17382 17724 17434
rect 17724 17382 17770 17434
rect 17474 17380 17530 17382
rect 17554 17380 17610 17382
rect 17634 17380 17690 17382
rect 17714 17380 17770 17382
rect 17474 16346 17530 16348
rect 17554 16346 17610 16348
rect 17634 16346 17690 16348
rect 17714 16346 17770 16348
rect 17474 16294 17520 16346
rect 17520 16294 17530 16346
rect 17554 16294 17584 16346
rect 17584 16294 17596 16346
rect 17596 16294 17610 16346
rect 17634 16294 17648 16346
rect 17648 16294 17660 16346
rect 17660 16294 17690 16346
rect 17714 16294 17724 16346
rect 17724 16294 17770 16346
rect 17474 16292 17530 16294
rect 17554 16292 17610 16294
rect 17634 16292 17690 16294
rect 17714 16292 17770 16294
rect 17474 15258 17530 15260
rect 17554 15258 17610 15260
rect 17634 15258 17690 15260
rect 17714 15258 17770 15260
rect 17474 15206 17520 15258
rect 17520 15206 17530 15258
rect 17554 15206 17584 15258
rect 17584 15206 17596 15258
rect 17596 15206 17610 15258
rect 17634 15206 17648 15258
rect 17648 15206 17660 15258
rect 17660 15206 17690 15258
rect 17714 15206 17724 15258
rect 17724 15206 17770 15258
rect 17474 15204 17530 15206
rect 17554 15204 17610 15206
rect 17634 15204 17690 15206
rect 17714 15204 17770 15206
rect 16814 13626 16870 13628
rect 16894 13626 16950 13628
rect 16974 13626 17030 13628
rect 17054 13626 17110 13628
rect 16814 13574 16860 13626
rect 16860 13574 16870 13626
rect 16894 13574 16924 13626
rect 16924 13574 16936 13626
rect 16936 13574 16950 13626
rect 16974 13574 16988 13626
rect 16988 13574 17000 13626
rect 17000 13574 17030 13626
rect 17054 13574 17064 13626
rect 17064 13574 17110 13626
rect 16814 13572 16870 13574
rect 16894 13572 16950 13574
rect 16974 13572 17030 13574
rect 17054 13572 17110 13574
rect 16814 12538 16870 12540
rect 16894 12538 16950 12540
rect 16974 12538 17030 12540
rect 17054 12538 17110 12540
rect 16814 12486 16860 12538
rect 16860 12486 16870 12538
rect 16894 12486 16924 12538
rect 16924 12486 16936 12538
rect 16936 12486 16950 12538
rect 16974 12486 16988 12538
rect 16988 12486 17000 12538
rect 17000 12486 17030 12538
rect 17054 12486 17064 12538
rect 17064 12486 17110 12538
rect 16814 12484 16870 12486
rect 16894 12484 16950 12486
rect 16974 12484 17030 12486
rect 17054 12484 17110 12486
rect 16814 11450 16870 11452
rect 16894 11450 16950 11452
rect 16974 11450 17030 11452
rect 17054 11450 17110 11452
rect 16814 11398 16860 11450
rect 16860 11398 16870 11450
rect 16894 11398 16924 11450
rect 16924 11398 16936 11450
rect 16936 11398 16950 11450
rect 16974 11398 16988 11450
rect 16988 11398 17000 11450
rect 17000 11398 17030 11450
rect 17054 11398 17064 11450
rect 17064 11398 17110 11450
rect 16814 11396 16870 11398
rect 16894 11396 16950 11398
rect 16974 11396 17030 11398
rect 17054 11396 17110 11398
rect 16814 10362 16870 10364
rect 16894 10362 16950 10364
rect 16974 10362 17030 10364
rect 17054 10362 17110 10364
rect 16814 10310 16860 10362
rect 16860 10310 16870 10362
rect 16894 10310 16924 10362
rect 16924 10310 16936 10362
rect 16936 10310 16950 10362
rect 16974 10310 16988 10362
rect 16988 10310 17000 10362
rect 17000 10310 17030 10362
rect 17054 10310 17064 10362
rect 17064 10310 17110 10362
rect 16814 10308 16870 10310
rect 16894 10308 16950 10310
rect 16974 10308 17030 10310
rect 17054 10308 17110 10310
rect 16814 9274 16870 9276
rect 16894 9274 16950 9276
rect 16974 9274 17030 9276
rect 17054 9274 17110 9276
rect 16814 9222 16860 9274
rect 16860 9222 16870 9274
rect 16894 9222 16924 9274
rect 16924 9222 16936 9274
rect 16936 9222 16950 9274
rect 16974 9222 16988 9274
rect 16988 9222 17000 9274
rect 17000 9222 17030 9274
rect 17054 9222 17064 9274
rect 17064 9222 17110 9274
rect 16814 9220 16870 9222
rect 16894 9220 16950 9222
rect 16974 9220 17030 9222
rect 17054 9220 17110 9222
rect 16814 8186 16870 8188
rect 16894 8186 16950 8188
rect 16974 8186 17030 8188
rect 17054 8186 17110 8188
rect 16814 8134 16860 8186
rect 16860 8134 16870 8186
rect 16894 8134 16924 8186
rect 16924 8134 16936 8186
rect 16936 8134 16950 8186
rect 16974 8134 16988 8186
rect 16988 8134 17000 8186
rect 17000 8134 17030 8186
rect 17054 8134 17064 8186
rect 17064 8134 17110 8186
rect 16814 8132 16870 8134
rect 16894 8132 16950 8134
rect 16974 8132 17030 8134
rect 17054 8132 17110 8134
rect 17474 14170 17530 14172
rect 17554 14170 17610 14172
rect 17634 14170 17690 14172
rect 17714 14170 17770 14172
rect 17474 14118 17520 14170
rect 17520 14118 17530 14170
rect 17554 14118 17584 14170
rect 17584 14118 17596 14170
rect 17596 14118 17610 14170
rect 17634 14118 17648 14170
rect 17648 14118 17660 14170
rect 17660 14118 17690 14170
rect 17714 14118 17724 14170
rect 17724 14118 17770 14170
rect 17474 14116 17530 14118
rect 17554 14116 17610 14118
rect 17634 14116 17690 14118
rect 17714 14116 17770 14118
rect 17474 13082 17530 13084
rect 17554 13082 17610 13084
rect 17634 13082 17690 13084
rect 17714 13082 17770 13084
rect 17474 13030 17520 13082
rect 17520 13030 17530 13082
rect 17554 13030 17584 13082
rect 17584 13030 17596 13082
rect 17596 13030 17610 13082
rect 17634 13030 17648 13082
rect 17648 13030 17660 13082
rect 17660 13030 17690 13082
rect 17714 13030 17724 13082
rect 17724 13030 17770 13082
rect 17474 13028 17530 13030
rect 17554 13028 17610 13030
rect 17634 13028 17690 13030
rect 17714 13028 17770 13030
rect 17474 11994 17530 11996
rect 17554 11994 17610 11996
rect 17634 11994 17690 11996
rect 17714 11994 17770 11996
rect 17474 11942 17520 11994
rect 17520 11942 17530 11994
rect 17554 11942 17584 11994
rect 17584 11942 17596 11994
rect 17596 11942 17610 11994
rect 17634 11942 17648 11994
rect 17648 11942 17660 11994
rect 17660 11942 17690 11994
rect 17714 11942 17724 11994
rect 17724 11942 17770 11994
rect 17474 11940 17530 11942
rect 17554 11940 17610 11942
rect 17634 11940 17690 11942
rect 17714 11940 17770 11942
rect 17474 10906 17530 10908
rect 17554 10906 17610 10908
rect 17634 10906 17690 10908
rect 17714 10906 17770 10908
rect 17474 10854 17520 10906
rect 17520 10854 17530 10906
rect 17554 10854 17584 10906
rect 17584 10854 17596 10906
rect 17596 10854 17610 10906
rect 17634 10854 17648 10906
rect 17648 10854 17660 10906
rect 17660 10854 17690 10906
rect 17714 10854 17724 10906
rect 17724 10854 17770 10906
rect 17474 10852 17530 10854
rect 17554 10852 17610 10854
rect 17634 10852 17690 10854
rect 17714 10852 17770 10854
rect 17474 9818 17530 9820
rect 17554 9818 17610 9820
rect 17634 9818 17690 9820
rect 17714 9818 17770 9820
rect 17474 9766 17520 9818
rect 17520 9766 17530 9818
rect 17554 9766 17584 9818
rect 17584 9766 17596 9818
rect 17596 9766 17610 9818
rect 17634 9766 17648 9818
rect 17648 9766 17660 9818
rect 17660 9766 17690 9818
rect 17714 9766 17724 9818
rect 17724 9766 17770 9818
rect 17474 9764 17530 9766
rect 17554 9764 17610 9766
rect 17634 9764 17690 9766
rect 17714 9764 17770 9766
rect 17474 8730 17530 8732
rect 17554 8730 17610 8732
rect 17634 8730 17690 8732
rect 17714 8730 17770 8732
rect 17474 8678 17520 8730
rect 17520 8678 17530 8730
rect 17554 8678 17584 8730
rect 17584 8678 17596 8730
rect 17596 8678 17610 8730
rect 17634 8678 17648 8730
rect 17648 8678 17660 8730
rect 17660 8678 17690 8730
rect 17714 8678 17724 8730
rect 17724 8678 17770 8730
rect 17474 8676 17530 8678
rect 17554 8676 17610 8678
rect 17634 8676 17690 8678
rect 17714 8676 17770 8678
rect 17474 7642 17530 7644
rect 17554 7642 17610 7644
rect 17634 7642 17690 7644
rect 17714 7642 17770 7644
rect 17474 7590 17520 7642
rect 17520 7590 17530 7642
rect 17554 7590 17584 7642
rect 17584 7590 17596 7642
rect 17596 7590 17610 7642
rect 17634 7590 17648 7642
rect 17648 7590 17660 7642
rect 17660 7590 17690 7642
rect 17714 7590 17724 7642
rect 17724 7590 17770 7642
rect 17474 7588 17530 7590
rect 17554 7588 17610 7590
rect 17634 7588 17690 7590
rect 17714 7588 17770 7590
rect 16814 7098 16870 7100
rect 16894 7098 16950 7100
rect 16974 7098 17030 7100
rect 17054 7098 17110 7100
rect 16814 7046 16860 7098
rect 16860 7046 16870 7098
rect 16894 7046 16924 7098
rect 16924 7046 16936 7098
rect 16936 7046 16950 7098
rect 16974 7046 16988 7098
rect 16988 7046 17000 7098
rect 17000 7046 17030 7098
rect 17054 7046 17064 7098
rect 17064 7046 17110 7098
rect 16814 7044 16870 7046
rect 16894 7044 16950 7046
rect 16974 7044 17030 7046
rect 17054 7044 17110 7046
rect 17474 6554 17530 6556
rect 17554 6554 17610 6556
rect 17634 6554 17690 6556
rect 17714 6554 17770 6556
rect 17474 6502 17520 6554
rect 17520 6502 17530 6554
rect 17554 6502 17584 6554
rect 17584 6502 17596 6554
rect 17596 6502 17610 6554
rect 17634 6502 17648 6554
rect 17648 6502 17660 6554
rect 17660 6502 17690 6554
rect 17714 6502 17724 6554
rect 17724 6502 17770 6554
rect 17474 6500 17530 6502
rect 17554 6500 17610 6502
rect 17634 6500 17690 6502
rect 17714 6500 17770 6502
rect 16814 6010 16870 6012
rect 16894 6010 16950 6012
rect 16974 6010 17030 6012
rect 17054 6010 17110 6012
rect 16814 5958 16860 6010
rect 16860 5958 16870 6010
rect 16894 5958 16924 6010
rect 16924 5958 16936 6010
rect 16936 5958 16950 6010
rect 16974 5958 16988 6010
rect 16988 5958 17000 6010
rect 17000 5958 17030 6010
rect 17054 5958 17064 6010
rect 17064 5958 17110 6010
rect 16814 5956 16870 5958
rect 16894 5956 16950 5958
rect 16974 5956 17030 5958
rect 17054 5956 17110 5958
rect 17474 5466 17530 5468
rect 17554 5466 17610 5468
rect 17634 5466 17690 5468
rect 17714 5466 17770 5468
rect 17474 5414 17520 5466
rect 17520 5414 17530 5466
rect 17554 5414 17584 5466
rect 17584 5414 17596 5466
rect 17596 5414 17610 5466
rect 17634 5414 17648 5466
rect 17648 5414 17660 5466
rect 17660 5414 17690 5466
rect 17714 5414 17724 5466
rect 17724 5414 17770 5466
rect 17474 5412 17530 5414
rect 17554 5412 17610 5414
rect 17634 5412 17690 5414
rect 17714 5412 17770 5414
rect 16814 4922 16870 4924
rect 16894 4922 16950 4924
rect 16974 4922 17030 4924
rect 17054 4922 17110 4924
rect 16814 4870 16860 4922
rect 16860 4870 16870 4922
rect 16894 4870 16924 4922
rect 16924 4870 16936 4922
rect 16936 4870 16950 4922
rect 16974 4870 16988 4922
rect 16988 4870 17000 4922
rect 17000 4870 17030 4922
rect 17054 4870 17064 4922
rect 17064 4870 17110 4922
rect 16814 4868 16870 4870
rect 16894 4868 16950 4870
rect 16974 4868 17030 4870
rect 17054 4868 17110 4870
rect 3881 4378 3937 4380
rect 3961 4378 4017 4380
rect 4041 4378 4097 4380
rect 4121 4378 4177 4380
rect 3881 4326 3927 4378
rect 3927 4326 3937 4378
rect 3961 4326 3991 4378
rect 3991 4326 4003 4378
rect 4003 4326 4017 4378
rect 4041 4326 4055 4378
rect 4055 4326 4067 4378
rect 4067 4326 4097 4378
rect 4121 4326 4131 4378
rect 4131 4326 4177 4378
rect 3881 4324 3937 4326
rect 3961 4324 4017 4326
rect 4041 4324 4097 4326
rect 4121 4324 4177 4326
rect 8412 4378 8468 4380
rect 8492 4378 8548 4380
rect 8572 4378 8628 4380
rect 8652 4378 8708 4380
rect 8412 4326 8458 4378
rect 8458 4326 8468 4378
rect 8492 4326 8522 4378
rect 8522 4326 8534 4378
rect 8534 4326 8548 4378
rect 8572 4326 8586 4378
rect 8586 4326 8598 4378
rect 8598 4326 8628 4378
rect 8652 4326 8662 4378
rect 8662 4326 8708 4378
rect 8412 4324 8468 4326
rect 8492 4324 8548 4326
rect 8572 4324 8628 4326
rect 8652 4324 8708 4326
rect 12943 4378 12999 4380
rect 13023 4378 13079 4380
rect 13103 4378 13159 4380
rect 13183 4378 13239 4380
rect 12943 4326 12989 4378
rect 12989 4326 12999 4378
rect 13023 4326 13053 4378
rect 13053 4326 13065 4378
rect 13065 4326 13079 4378
rect 13103 4326 13117 4378
rect 13117 4326 13129 4378
rect 13129 4326 13159 4378
rect 13183 4326 13193 4378
rect 13193 4326 13239 4378
rect 12943 4324 12999 4326
rect 13023 4324 13079 4326
rect 13103 4324 13159 4326
rect 13183 4324 13239 4326
rect 17474 4378 17530 4380
rect 17554 4378 17610 4380
rect 17634 4378 17690 4380
rect 17714 4378 17770 4380
rect 17474 4326 17520 4378
rect 17520 4326 17530 4378
rect 17554 4326 17584 4378
rect 17584 4326 17596 4378
rect 17596 4326 17610 4378
rect 17634 4326 17648 4378
rect 17648 4326 17660 4378
rect 17660 4326 17690 4378
rect 17714 4326 17724 4378
rect 17724 4326 17770 4378
rect 17474 4324 17530 4326
rect 17554 4324 17610 4326
rect 17634 4324 17690 4326
rect 17714 4324 17770 4326
rect 3221 3834 3277 3836
rect 3301 3834 3357 3836
rect 3381 3834 3437 3836
rect 3461 3834 3517 3836
rect 3221 3782 3267 3834
rect 3267 3782 3277 3834
rect 3301 3782 3331 3834
rect 3331 3782 3343 3834
rect 3343 3782 3357 3834
rect 3381 3782 3395 3834
rect 3395 3782 3407 3834
rect 3407 3782 3437 3834
rect 3461 3782 3471 3834
rect 3471 3782 3517 3834
rect 3221 3780 3277 3782
rect 3301 3780 3357 3782
rect 3381 3780 3437 3782
rect 3461 3780 3517 3782
rect 7752 3834 7808 3836
rect 7832 3834 7888 3836
rect 7912 3834 7968 3836
rect 7992 3834 8048 3836
rect 7752 3782 7798 3834
rect 7798 3782 7808 3834
rect 7832 3782 7862 3834
rect 7862 3782 7874 3834
rect 7874 3782 7888 3834
rect 7912 3782 7926 3834
rect 7926 3782 7938 3834
rect 7938 3782 7968 3834
rect 7992 3782 8002 3834
rect 8002 3782 8048 3834
rect 7752 3780 7808 3782
rect 7832 3780 7888 3782
rect 7912 3780 7968 3782
rect 7992 3780 8048 3782
rect 12283 3834 12339 3836
rect 12363 3834 12419 3836
rect 12443 3834 12499 3836
rect 12523 3834 12579 3836
rect 12283 3782 12329 3834
rect 12329 3782 12339 3834
rect 12363 3782 12393 3834
rect 12393 3782 12405 3834
rect 12405 3782 12419 3834
rect 12443 3782 12457 3834
rect 12457 3782 12469 3834
rect 12469 3782 12499 3834
rect 12523 3782 12533 3834
rect 12533 3782 12579 3834
rect 12283 3780 12339 3782
rect 12363 3780 12419 3782
rect 12443 3780 12499 3782
rect 12523 3780 12579 3782
rect 3881 3290 3937 3292
rect 3961 3290 4017 3292
rect 4041 3290 4097 3292
rect 4121 3290 4177 3292
rect 3881 3238 3927 3290
rect 3927 3238 3937 3290
rect 3961 3238 3991 3290
rect 3991 3238 4003 3290
rect 4003 3238 4017 3290
rect 4041 3238 4055 3290
rect 4055 3238 4067 3290
rect 4067 3238 4097 3290
rect 4121 3238 4131 3290
rect 4131 3238 4177 3290
rect 3881 3236 3937 3238
rect 3961 3236 4017 3238
rect 4041 3236 4097 3238
rect 4121 3236 4177 3238
rect 8412 3290 8468 3292
rect 8492 3290 8548 3292
rect 8572 3290 8628 3292
rect 8652 3290 8708 3292
rect 8412 3238 8458 3290
rect 8458 3238 8468 3290
rect 8492 3238 8522 3290
rect 8522 3238 8534 3290
rect 8534 3238 8548 3290
rect 8572 3238 8586 3290
rect 8586 3238 8598 3290
rect 8598 3238 8628 3290
rect 8652 3238 8662 3290
rect 8662 3238 8708 3290
rect 8412 3236 8468 3238
rect 8492 3236 8548 3238
rect 8572 3236 8628 3238
rect 8652 3236 8708 3238
rect 12943 3290 12999 3292
rect 13023 3290 13079 3292
rect 13103 3290 13159 3292
rect 13183 3290 13239 3292
rect 12943 3238 12989 3290
rect 12989 3238 12999 3290
rect 13023 3238 13053 3290
rect 13053 3238 13065 3290
rect 13065 3238 13079 3290
rect 13103 3238 13117 3290
rect 13117 3238 13129 3290
rect 13129 3238 13159 3290
rect 13183 3238 13193 3290
rect 13193 3238 13239 3290
rect 12943 3236 12999 3238
rect 13023 3236 13079 3238
rect 13103 3236 13159 3238
rect 13183 3236 13239 3238
rect 3221 2746 3277 2748
rect 3301 2746 3357 2748
rect 3381 2746 3437 2748
rect 3461 2746 3517 2748
rect 3221 2694 3267 2746
rect 3267 2694 3277 2746
rect 3301 2694 3331 2746
rect 3331 2694 3343 2746
rect 3343 2694 3357 2746
rect 3381 2694 3395 2746
rect 3395 2694 3407 2746
rect 3407 2694 3437 2746
rect 3461 2694 3471 2746
rect 3471 2694 3517 2746
rect 3221 2692 3277 2694
rect 3301 2692 3357 2694
rect 3381 2692 3437 2694
rect 3461 2692 3517 2694
rect 7752 2746 7808 2748
rect 7832 2746 7888 2748
rect 7912 2746 7968 2748
rect 7992 2746 8048 2748
rect 7752 2694 7798 2746
rect 7798 2694 7808 2746
rect 7832 2694 7862 2746
rect 7862 2694 7874 2746
rect 7874 2694 7888 2746
rect 7912 2694 7926 2746
rect 7926 2694 7938 2746
rect 7938 2694 7968 2746
rect 7992 2694 8002 2746
rect 8002 2694 8048 2746
rect 7752 2692 7808 2694
rect 7832 2692 7888 2694
rect 7912 2692 7968 2694
rect 7992 2692 8048 2694
rect 12283 2746 12339 2748
rect 12363 2746 12419 2748
rect 12443 2746 12499 2748
rect 12523 2746 12579 2748
rect 12283 2694 12329 2746
rect 12329 2694 12339 2746
rect 12363 2694 12393 2746
rect 12393 2694 12405 2746
rect 12405 2694 12419 2746
rect 12443 2694 12457 2746
rect 12457 2694 12469 2746
rect 12469 2694 12499 2746
rect 12523 2694 12533 2746
rect 12533 2694 12579 2746
rect 12283 2692 12339 2694
rect 12363 2692 12419 2694
rect 12443 2692 12499 2694
rect 12523 2692 12579 2694
rect 16814 3834 16870 3836
rect 16894 3834 16950 3836
rect 16974 3834 17030 3836
rect 17054 3834 17110 3836
rect 16814 3782 16860 3834
rect 16860 3782 16870 3834
rect 16894 3782 16924 3834
rect 16924 3782 16936 3834
rect 16936 3782 16950 3834
rect 16974 3782 16988 3834
rect 16988 3782 17000 3834
rect 17000 3782 17030 3834
rect 17054 3782 17064 3834
rect 17064 3782 17110 3834
rect 16814 3780 16870 3782
rect 16894 3780 16950 3782
rect 16974 3780 17030 3782
rect 17054 3780 17110 3782
rect 17474 3290 17530 3292
rect 17554 3290 17610 3292
rect 17634 3290 17690 3292
rect 17714 3290 17770 3292
rect 17474 3238 17520 3290
rect 17520 3238 17530 3290
rect 17554 3238 17584 3290
rect 17584 3238 17596 3290
rect 17596 3238 17610 3290
rect 17634 3238 17648 3290
rect 17648 3238 17660 3290
rect 17660 3238 17690 3290
rect 17714 3238 17724 3290
rect 17724 3238 17770 3290
rect 17474 3236 17530 3238
rect 17554 3236 17610 3238
rect 17634 3236 17690 3238
rect 17714 3236 17770 3238
rect 16814 2746 16870 2748
rect 16894 2746 16950 2748
rect 16974 2746 17030 2748
rect 17054 2746 17110 2748
rect 16814 2694 16860 2746
rect 16860 2694 16870 2746
rect 16894 2694 16924 2746
rect 16924 2694 16936 2746
rect 16936 2694 16950 2746
rect 16974 2694 16988 2746
rect 16988 2694 17000 2746
rect 17000 2694 17030 2746
rect 17054 2694 17064 2746
rect 17064 2694 17110 2746
rect 16814 2692 16870 2694
rect 16894 2692 16950 2694
rect 16974 2692 17030 2694
rect 17054 2692 17110 2694
rect 3881 2202 3937 2204
rect 3961 2202 4017 2204
rect 4041 2202 4097 2204
rect 4121 2202 4177 2204
rect 3881 2150 3927 2202
rect 3927 2150 3937 2202
rect 3961 2150 3991 2202
rect 3991 2150 4003 2202
rect 4003 2150 4017 2202
rect 4041 2150 4055 2202
rect 4055 2150 4067 2202
rect 4067 2150 4097 2202
rect 4121 2150 4131 2202
rect 4131 2150 4177 2202
rect 3881 2148 3937 2150
rect 3961 2148 4017 2150
rect 4041 2148 4097 2150
rect 4121 2148 4177 2150
rect 8412 2202 8468 2204
rect 8492 2202 8548 2204
rect 8572 2202 8628 2204
rect 8652 2202 8708 2204
rect 8412 2150 8458 2202
rect 8458 2150 8468 2202
rect 8492 2150 8522 2202
rect 8522 2150 8534 2202
rect 8534 2150 8548 2202
rect 8572 2150 8586 2202
rect 8586 2150 8598 2202
rect 8598 2150 8628 2202
rect 8652 2150 8662 2202
rect 8662 2150 8708 2202
rect 8412 2148 8468 2150
rect 8492 2148 8548 2150
rect 8572 2148 8628 2150
rect 8652 2148 8708 2150
rect 12943 2202 12999 2204
rect 13023 2202 13079 2204
rect 13103 2202 13159 2204
rect 13183 2202 13239 2204
rect 12943 2150 12989 2202
rect 12989 2150 12999 2202
rect 13023 2150 13053 2202
rect 13053 2150 13065 2202
rect 13065 2150 13079 2202
rect 13103 2150 13117 2202
rect 13117 2150 13129 2202
rect 13129 2150 13159 2202
rect 13183 2150 13193 2202
rect 13193 2150 13239 2202
rect 12943 2148 12999 2150
rect 13023 2148 13079 2150
rect 13103 2148 13159 2150
rect 13183 2148 13239 2150
rect 17474 2202 17530 2204
rect 17554 2202 17610 2204
rect 17634 2202 17690 2204
rect 17714 2202 17770 2204
rect 17474 2150 17520 2202
rect 17520 2150 17530 2202
rect 17554 2150 17584 2202
rect 17584 2150 17596 2202
rect 17596 2150 17610 2202
rect 17634 2150 17648 2202
rect 17648 2150 17660 2202
rect 17660 2150 17690 2202
rect 17714 2150 17724 2202
rect 17724 2150 17770 2202
rect 17474 2148 17530 2150
rect 17554 2148 17610 2150
rect 17634 2148 17690 2150
rect 17714 2148 17770 2150
<< metal3 >>
rect 3211 20160 3527 20161
rect 3211 20096 3217 20160
rect 3281 20096 3297 20160
rect 3361 20096 3377 20160
rect 3441 20096 3457 20160
rect 3521 20096 3527 20160
rect 3211 20095 3527 20096
rect 7742 20160 8058 20161
rect 7742 20096 7748 20160
rect 7812 20096 7828 20160
rect 7892 20096 7908 20160
rect 7972 20096 7988 20160
rect 8052 20096 8058 20160
rect 7742 20095 8058 20096
rect 12273 20160 12589 20161
rect 12273 20096 12279 20160
rect 12343 20096 12359 20160
rect 12423 20096 12439 20160
rect 12503 20096 12519 20160
rect 12583 20096 12589 20160
rect 12273 20095 12589 20096
rect 16804 20160 17120 20161
rect 16804 20096 16810 20160
rect 16874 20096 16890 20160
rect 16954 20096 16970 20160
rect 17034 20096 17050 20160
rect 17114 20096 17120 20160
rect 16804 20095 17120 20096
rect 17125 19818 17191 19821
rect 17677 19818 17743 19821
rect 17125 19816 17743 19818
rect 17125 19760 17130 19816
rect 17186 19760 17682 19816
rect 17738 19760 17743 19816
rect 17125 19758 17743 19760
rect 17125 19755 17191 19758
rect 17677 19755 17743 19758
rect 3871 19616 4187 19617
rect 3871 19552 3877 19616
rect 3941 19552 3957 19616
rect 4021 19552 4037 19616
rect 4101 19552 4117 19616
rect 4181 19552 4187 19616
rect 3871 19551 4187 19552
rect 8402 19616 8718 19617
rect 8402 19552 8408 19616
rect 8472 19552 8488 19616
rect 8552 19552 8568 19616
rect 8632 19552 8648 19616
rect 8712 19552 8718 19616
rect 8402 19551 8718 19552
rect 12933 19616 13249 19617
rect 12933 19552 12939 19616
rect 13003 19552 13019 19616
rect 13083 19552 13099 19616
rect 13163 19552 13179 19616
rect 13243 19552 13249 19616
rect 12933 19551 13249 19552
rect 17464 19616 17780 19617
rect 17464 19552 17470 19616
rect 17534 19552 17550 19616
rect 17614 19552 17630 19616
rect 17694 19552 17710 19616
rect 17774 19552 17780 19616
rect 17464 19551 17780 19552
rect 3211 19072 3527 19073
rect 3211 19008 3217 19072
rect 3281 19008 3297 19072
rect 3361 19008 3377 19072
rect 3441 19008 3457 19072
rect 3521 19008 3527 19072
rect 3211 19007 3527 19008
rect 7742 19072 8058 19073
rect 7742 19008 7748 19072
rect 7812 19008 7828 19072
rect 7892 19008 7908 19072
rect 7972 19008 7988 19072
rect 8052 19008 8058 19072
rect 7742 19007 8058 19008
rect 12273 19072 12589 19073
rect 12273 19008 12279 19072
rect 12343 19008 12359 19072
rect 12423 19008 12439 19072
rect 12503 19008 12519 19072
rect 12583 19008 12589 19072
rect 12273 19007 12589 19008
rect 16804 19072 17120 19073
rect 16804 19008 16810 19072
rect 16874 19008 16890 19072
rect 16954 19008 16970 19072
rect 17034 19008 17050 19072
rect 17114 19008 17120 19072
rect 16804 19007 17120 19008
rect 3871 18528 4187 18529
rect 3871 18464 3877 18528
rect 3941 18464 3957 18528
rect 4021 18464 4037 18528
rect 4101 18464 4117 18528
rect 4181 18464 4187 18528
rect 3871 18463 4187 18464
rect 8402 18528 8718 18529
rect 8402 18464 8408 18528
rect 8472 18464 8488 18528
rect 8552 18464 8568 18528
rect 8632 18464 8648 18528
rect 8712 18464 8718 18528
rect 8402 18463 8718 18464
rect 12933 18528 13249 18529
rect 12933 18464 12939 18528
rect 13003 18464 13019 18528
rect 13083 18464 13099 18528
rect 13163 18464 13179 18528
rect 13243 18464 13249 18528
rect 12933 18463 13249 18464
rect 17464 18528 17780 18529
rect 17464 18464 17470 18528
rect 17534 18464 17550 18528
rect 17614 18464 17630 18528
rect 17694 18464 17710 18528
rect 17774 18464 17780 18528
rect 17464 18463 17780 18464
rect 3211 17984 3527 17985
rect 3211 17920 3217 17984
rect 3281 17920 3297 17984
rect 3361 17920 3377 17984
rect 3441 17920 3457 17984
rect 3521 17920 3527 17984
rect 3211 17919 3527 17920
rect 7742 17984 8058 17985
rect 7742 17920 7748 17984
rect 7812 17920 7828 17984
rect 7892 17920 7908 17984
rect 7972 17920 7988 17984
rect 8052 17920 8058 17984
rect 7742 17919 8058 17920
rect 12273 17984 12589 17985
rect 12273 17920 12279 17984
rect 12343 17920 12359 17984
rect 12423 17920 12439 17984
rect 12503 17920 12519 17984
rect 12583 17920 12589 17984
rect 12273 17919 12589 17920
rect 16804 17984 17120 17985
rect 16804 17920 16810 17984
rect 16874 17920 16890 17984
rect 16954 17920 16970 17984
rect 17034 17920 17050 17984
rect 17114 17920 17120 17984
rect 16804 17919 17120 17920
rect 3871 17440 4187 17441
rect 3871 17376 3877 17440
rect 3941 17376 3957 17440
rect 4021 17376 4037 17440
rect 4101 17376 4117 17440
rect 4181 17376 4187 17440
rect 3871 17375 4187 17376
rect 8402 17440 8718 17441
rect 8402 17376 8408 17440
rect 8472 17376 8488 17440
rect 8552 17376 8568 17440
rect 8632 17376 8648 17440
rect 8712 17376 8718 17440
rect 8402 17375 8718 17376
rect 12933 17440 13249 17441
rect 12933 17376 12939 17440
rect 13003 17376 13019 17440
rect 13083 17376 13099 17440
rect 13163 17376 13179 17440
rect 13243 17376 13249 17440
rect 12933 17375 13249 17376
rect 17464 17440 17780 17441
rect 17464 17376 17470 17440
rect 17534 17376 17550 17440
rect 17614 17376 17630 17440
rect 17694 17376 17710 17440
rect 17774 17376 17780 17440
rect 17464 17375 17780 17376
rect 3211 16896 3527 16897
rect 3211 16832 3217 16896
rect 3281 16832 3297 16896
rect 3361 16832 3377 16896
rect 3441 16832 3457 16896
rect 3521 16832 3527 16896
rect 3211 16831 3527 16832
rect 7742 16896 8058 16897
rect 7742 16832 7748 16896
rect 7812 16832 7828 16896
rect 7892 16832 7908 16896
rect 7972 16832 7988 16896
rect 8052 16832 8058 16896
rect 7742 16831 8058 16832
rect 12273 16896 12589 16897
rect 12273 16832 12279 16896
rect 12343 16832 12359 16896
rect 12423 16832 12439 16896
rect 12503 16832 12519 16896
rect 12583 16832 12589 16896
rect 12273 16831 12589 16832
rect 16804 16896 17120 16897
rect 16804 16832 16810 16896
rect 16874 16832 16890 16896
rect 16954 16832 16970 16896
rect 17034 16832 17050 16896
rect 17114 16832 17120 16896
rect 16804 16831 17120 16832
rect 0 16690 800 16720
rect 933 16690 999 16693
rect 0 16688 999 16690
rect 0 16632 938 16688
rect 994 16632 999 16688
rect 0 16630 999 16632
rect 0 16600 800 16630
rect 933 16627 999 16630
rect 3871 16352 4187 16353
rect 3871 16288 3877 16352
rect 3941 16288 3957 16352
rect 4021 16288 4037 16352
rect 4101 16288 4117 16352
rect 4181 16288 4187 16352
rect 3871 16287 4187 16288
rect 8402 16352 8718 16353
rect 8402 16288 8408 16352
rect 8472 16288 8488 16352
rect 8552 16288 8568 16352
rect 8632 16288 8648 16352
rect 8712 16288 8718 16352
rect 8402 16287 8718 16288
rect 12933 16352 13249 16353
rect 12933 16288 12939 16352
rect 13003 16288 13019 16352
rect 13083 16288 13099 16352
rect 13163 16288 13179 16352
rect 13243 16288 13249 16352
rect 12933 16287 13249 16288
rect 17464 16352 17780 16353
rect 17464 16288 17470 16352
rect 17534 16288 17550 16352
rect 17614 16288 17630 16352
rect 17694 16288 17710 16352
rect 17774 16288 17780 16352
rect 17464 16287 17780 16288
rect 3211 15808 3527 15809
rect 3211 15744 3217 15808
rect 3281 15744 3297 15808
rect 3361 15744 3377 15808
rect 3441 15744 3457 15808
rect 3521 15744 3527 15808
rect 3211 15743 3527 15744
rect 7742 15808 8058 15809
rect 7742 15744 7748 15808
rect 7812 15744 7828 15808
rect 7892 15744 7908 15808
rect 7972 15744 7988 15808
rect 8052 15744 8058 15808
rect 7742 15743 8058 15744
rect 12273 15808 12589 15809
rect 12273 15744 12279 15808
rect 12343 15744 12359 15808
rect 12423 15744 12439 15808
rect 12503 15744 12519 15808
rect 12583 15744 12589 15808
rect 12273 15743 12589 15744
rect 16804 15808 17120 15809
rect 16804 15744 16810 15808
rect 16874 15744 16890 15808
rect 16954 15744 16970 15808
rect 17034 15744 17050 15808
rect 17114 15744 17120 15808
rect 16804 15743 17120 15744
rect 3871 15264 4187 15265
rect 3871 15200 3877 15264
rect 3941 15200 3957 15264
rect 4021 15200 4037 15264
rect 4101 15200 4117 15264
rect 4181 15200 4187 15264
rect 3871 15199 4187 15200
rect 8402 15264 8718 15265
rect 8402 15200 8408 15264
rect 8472 15200 8488 15264
rect 8552 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8718 15264
rect 8402 15199 8718 15200
rect 12933 15264 13249 15265
rect 12933 15200 12939 15264
rect 13003 15200 13019 15264
rect 13083 15200 13099 15264
rect 13163 15200 13179 15264
rect 13243 15200 13249 15264
rect 12933 15199 13249 15200
rect 17464 15264 17780 15265
rect 17464 15200 17470 15264
rect 17534 15200 17550 15264
rect 17614 15200 17630 15264
rect 17694 15200 17710 15264
rect 17774 15200 17780 15264
rect 17464 15199 17780 15200
rect 3211 14720 3527 14721
rect 3211 14656 3217 14720
rect 3281 14656 3297 14720
rect 3361 14656 3377 14720
rect 3441 14656 3457 14720
rect 3521 14656 3527 14720
rect 3211 14655 3527 14656
rect 7742 14720 8058 14721
rect 7742 14656 7748 14720
rect 7812 14656 7828 14720
rect 7892 14656 7908 14720
rect 7972 14656 7988 14720
rect 8052 14656 8058 14720
rect 7742 14655 8058 14656
rect 12273 14720 12589 14721
rect 12273 14656 12279 14720
rect 12343 14656 12359 14720
rect 12423 14656 12439 14720
rect 12503 14656 12519 14720
rect 12583 14656 12589 14720
rect 12273 14655 12589 14656
rect 16804 14720 17120 14721
rect 16804 14656 16810 14720
rect 16874 14656 16890 14720
rect 16954 14656 16970 14720
rect 17034 14656 17050 14720
rect 17114 14656 17120 14720
rect 16804 14655 17120 14656
rect 3871 14176 4187 14177
rect 3871 14112 3877 14176
rect 3941 14112 3957 14176
rect 4021 14112 4037 14176
rect 4101 14112 4117 14176
rect 4181 14112 4187 14176
rect 3871 14111 4187 14112
rect 8402 14176 8718 14177
rect 8402 14112 8408 14176
rect 8472 14112 8488 14176
rect 8552 14112 8568 14176
rect 8632 14112 8648 14176
rect 8712 14112 8718 14176
rect 8402 14111 8718 14112
rect 12933 14176 13249 14177
rect 12933 14112 12939 14176
rect 13003 14112 13019 14176
rect 13083 14112 13099 14176
rect 13163 14112 13179 14176
rect 13243 14112 13249 14176
rect 12933 14111 13249 14112
rect 17464 14176 17780 14177
rect 17464 14112 17470 14176
rect 17534 14112 17550 14176
rect 17614 14112 17630 14176
rect 17694 14112 17710 14176
rect 17774 14112 17780 14176
rect 17464 14111 17780 14112
rect 3211 13632 3527 13633
rect 3211 13568 3217 13632
rect 3281 13568 3297 13632
rect 3361 13568 3377 13632
rect 3441 13568 3457 13632
rect 3521 13568 3527 13632
rect 3211 13567 3527 13568
rect 7742 13632 8058 13633
rect 7742 13568 7748 13632
rect 7812 13568 7828 13632
rect 7892 13568 7908 13632
rect 7972 13568 7988 13632
rect 8052 13568 8058 13632
rect 7742 13567 8058 13568
rect 12273 13632 12589 13633
rect 12273 13568 12279 13632
rect 12343 13568 12359 13632
rect 12423 13568 12439 13632
rect 12503 13568 12519 13632
rect 12583 13568 12589 13632
rect 12273 13567 12589 13568
rect 16804 13632 17120 13633
rect 16804 13568 16810 13632
rect 16874 13568 16890 13632
rect 16954 13568 16970 13632
rect 17034 13568 17050 13632
rect 17114 13568 17120 13632
rect 16804 13567 17120 13568
rect 3871 13088 4187 13089
rect 3871 13024 3877 13088
rect 3941 13024 3957 13088
rect 4021 13024 4037 13088
rect 4101 13024 4117 13088
rect 4181 13024 4187 13088
rect 3871 13023 4187 13024
rect 8402 13088 8718 13089
rect 8402 13024 8408 13088
rect 8472 13024 8488 13088
rect 8552 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8718 13088
rect 8402 13023 8718 13024
rect 12933 13088 13249 13089
rect 12933 13024 12939 13088
rect 13003 13024 13019 13088
rect 13083 13024 13099 13088
rect 13163 13024 13179 13088
rect 13243 13024 13249 13088
rect 12933 13023 13249 13024
rect 17464 13088 17780 13089
rect 17464 13024 17470 13088
rect 17534 13024 17550 13088
rect 17614 13024 17630 13088
rect 17694 13024 17710 13088
rect 17774 13024 17780 13088
rect 17464 13023 17780 13024
rect 2681 12882 2747 12885
rect 2681 12880 4354 12882
rect 2681 12824 2686 12880
rect 2742 12824 4354 12880
rect 2681 12822 4354 12824
rect 2681 12819 2747 12822
rect 3211 12544 3527 12545
rect 3211 12480 3217 12544
rect 3281 12480 3297 12544
rect 3361 12480 3377 12544
rect 3441 12480 3457 12544
rect 3521 12480 3527 12544
rect 3211 12479 3527 12480
rect 4294 12476 4354 12822
rect 7742 12544 8058 12545
rect 7742 12480 7748 12544
rect 7812 12480 7828 12544
rect 7892 12480 7908 12544
rect 7972 12480 7988 12544
rect 8052 12480 8058 12544
rect 7742 12479 8058 12480
rect 12273 12544 12589 12545
rect 12273 12480 12279 12544
rect 12343 12480 12359 12544
rect 12423 12480 12439 12544
rect 12503 12480 12519 12544
rect 12583 12480 12589 12544
rect 12273 12479 12589 12480
rect 16804 12544 17120 12545
rect 16804 12480 16810 12544
rect 16874 12480 16890 12544
rect 16954 12480 16970 12544
rect 17034 12480 17050 12544
rect 17114 12480 17120 12544
rect 16804 12479 17120 12480
rect 4286 12412 4292 12476
rect 4356 12474 4362 12476
rect 5257 12474 5323 12477
rect 4356 12472 5323 12474
rect 4356 12416 5262 12472
rect 5318 12416 5323 12472
rect 4356 12414 5323 12416
rect 4356 12412 4362 12414
rect 5257 12411 5323 12414
rect 5257 12338 5323 12341
rect 9765 12338 9831 12341
rect 12801 12338 12867 12341
rect 5257 12336 12867 12338
rect 5257 12280 5262 12336
rect 5318 12280 9770 12336
rect 9826 12280 12806 12336
rect 12862 12280 12867 12336
rect 5257 12278 12867 12280
rect 5257 12275 5323 12278
rect 9765 12275 9831 12278
rect 12801 12275 12867 12278
rect 3871 12000 4187 12001
rect 3871 11936 3877 12000
rect 3941 11936 3957 12000
rect 4021 11936 4037 12000
rect 4101 11936 4117 12000
rect 4181 11936 4187 12000
rect 3871 11935 4187 11936
rect 8402 12000 8718 12001
rect 8402 11936 8408 12000
rect 8472 11936 8488 12000
rect 8552 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8718 12000
rect 8402 11935 8718 11936
rect 12933 12000 13249 12001
rect 12933 11936 12939 12000
rect 13003 11936 13019 12000
rect 13083 11936 13099 12000
rect 13163 11936 13179 12000
rect 13243 11936 13249 12000
rect 12933 11935 13249 11936
rect 17464 12000 17780 12001
rect 17464 11936 17470 12000
rect 17534 11936 17550 12000
rect 17614 11936 17630 12000
rect 17694 11936 17710 12000
rect 17774 11936 17780 12000
rect 17464 11935 17780 11936
rect 3211 11456 3527 11457
rect 3211 11392 3217 11456
rect 3281 11392 3297 11456
rect 3361 11392 3377 11456
rect 3441 11392 3457 11456
rect 3521 11392 3527 11456
rect 3211 11391 3527 11392
rect 7742 11456 8058 11457
rect 7742 11392 7748 11456
rect 7812 11392 7828 11456
rect 7892 11392 7908 11456
rect 7972 11392 7988 11456
rect 8052 11392 8058 11456
rect 7742 11391 8058 11392
rect 12273 11456 12589 11457
rect 12273 11392 12279 11456
rect 12343 11392 12359 11456
rect 12423 11392 12439 11456
rect 12503 11392 12519 11456
rect 12583 11392 12589 11456
rect 12273 11391 12589 11392
rect 16804 11456 17120 11457
rect 16804 11392 16810 11456
rect 16874 11392 16890 11456
rect 16954 11392 16970 11456
rect 17034 11392 17050 11456
rect 17114 11392 17120 11456
rect 16804 11391 17120 11392
rect 11053 11250 11119 11253
rect 19570 11250 20370 11280
rect 11053 11248 20370 11250
rect 11053 11192 11058 11248
rect 11114 11192 20370 11248
rect 11053 11190 20370 11192
rect 11053 11187 11119 11190
rect 19570 11160 20370 11190
rect 3871 10912 4187 10913
rect 3871 10848 3877 10912
rect 3941 10848 3957 10912
rect 4021 10848 4037 10912
rect 4101 10848 4117 10912
rect 4181 10848 4187 10912
rect 3871 10847 4187 10848
rect 8402 10912 8718 10913
rect 8402 10848 8408 10912
rect 8472 10848 8488 10912
rect 8552 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8718 10912
rect 8402 10847 8718 10848
rect 12933 10912 13249 10913
rect 12933 10848 12939 10912
rect 13003 10848 13019 10912
rect 13083 10848 13099 10912
rect 13163 10848 13179 10912
rect 13243 10848 13249 10912
rect 12933 10847 13249 10848
rect 17464 10912 17780 10913
rect 17464 10848 17470 10912
rect 17534 10848 17550 10912
rect 17614 10848 17630 10912
rect 17694 10848 17710 10912
rect 17774 10848 17780 10912
rect 17464 10847 17780 10848
rect 3211 10368 3527 10369
rect 3211 10304 3217 10368
rect 3281 10304 3297 10368
rect 3361 10304 3377 10368
rect 3441 10304 3457 10368
rect 3521 10304 3527 10368
rect 3211 10303 3527 10304
rect 7742 10368 8058 10369
rect 7742 10304 7748 10368
rect 7812 10304 7828 10368
rect 7892 10304 7908 10368
rect 7972 10304 7988 10368
rect 8052 10304 8058 10368
rect 7742 10303 8058 10304
rect 12273 10368 12589 10369
rect 12273 10304 12279 10368
rect 12343 10304 12359 10368
rect 12423 10304 12439 10368
rect 12503 10304 12519 10368
rect 12583 10304 12589 10368
rect 12273 10303 12589 10304
rect 16804 10368 17120 10369
rect 16804 10304 16810 10368
rect 16874 10304 16890 10368
rect 16954 10304 16970 10368
rect 17034 10304 17050 10368
rect 17114 10304 17120 10368
rect 16804 10303 17120 10304
rect 3871 9824 4187 9825
rect 3871 9760 3877 9824
rect 3941 9760 3957 9824
rect 4021 9760 4037 9824
rect 4101 9760 4117 9824
rect 4181 9760 4187 9824
rect 3871 9759 4187 9760
rect 8402 9824 8718 9825
rect 8402 9760 8408 9824
rect 8472 9760 8488 9824
rect 8552 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8718 9824
rect 8402 9759 8718 9760
rect 12933 9824 13249 9825
rect 12933 9760 12939 9824
rect 13003 9760 13019 9824
rect 13083 9760 13099 9824
rect 13163 9760 13179 9824
rect 13243 9760 13249 9824
rect 12933 9759 13249 9760
rect 17464 9824 17780 9825
rect 17464 9760 17470 9824
rect 17534 9760 17550 9824
rect 17614 9760 17630 9824
rect 17694 9760 17710 9824
rect 17774 9760 17780 9824
rect 17464 9759 17780 9760
rect 3211 9280 3527 9281
rect 3211 9216 3217 9280
rect 3281 9216 3297 9280
rect 3361 9216 3377 9280
rect 3441 9216 3457 9280
rect 3521 9216 3527 9280
rect 3211 9215 3527 9216
rect 7742 9280 8058 9281
rect 7742 9216 7748 9280
rect 7812 9216 7828 9280
rect 7892 9216 7908 9280
rect 7972 9216 7988 9280
rect 8052 9216 8058 9280
rect 7742 9215 8058 9216
rect 12273 9280 12589 9281
rect 12273 9216 12279 9280
rect 12343 9216 12359 9280
rect 12423 9216 12439 9280
rect 12503 9216 12519 9280
rect 12583 9216 12589 9280
rect 12273 9215 12589 9216
rect 16804 9280 17120 9281
rect 16804 9216 16810 9280
rect 16874 9216 16890 9280
rect 16954 9216 16970 9280
rect 17034 9216 17050 9280
rect 17114 9216 17120 9280
rect 16804 9215 17120 9216
rect 3871 8736 4187 8737
rect 3871 8672 3877 8736
rect 3941 8672 3957 8736
rect 4021 8672 4037 8736
rect 4101 8672 4117 8736
rect 4181 8672 4187 8736
rect 3871 8671 4187 8672
rect 8402 8736 8718 8737
rect 8402 8672 8408 8736
rect 8472 8672 8488 8736
rect 8552 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8718 8736
rect 8402 8671 8718 8672
rect 12933 8736 13249 8737
rect 12933 8672 12939 8736
rect 13003 8672 13019 8736
rect 13083 8672 13099 8736
rect 13163 8672 13179 8736
rect 13243 8672 13249 8736
rect 12933 8671 13249 8672
rect 17464 8736 17780 8737
rect 17464 8672 17470 8736
rect 17534 8672 17550 8736
rect 17614 8672 17630 8736
rect 17694 8672 17710 8736
rect 17774 8672 17780 8736
rect 17464 8671 17780 8672
rect 4153 8258 4219 8261
rect 4286 8258 4292 8260
rect 4153 8256 4292 8258
rect 4153 8200 4158 8256
rect 4214 8200 4292 8256
rect 4153 8198 4292 8200
rect 4153 8195 4219 8198
rect 4286 8196 4292 8198
rect 4356 8196 4362 8260
rect 3211 8192 3527 8193
rect 3211 8128 3217 8192
rect 3281 8128 3297 8192
rect 3361 8128 3377 8192
rect 3441 8128 3457 8192
rect 3521 8128 3527 8192
rect 3211 8127 3527 8128
rect 7742 8192 8058 8193
rect 7742 8128 7748 8192
rect 7812 8128 7828 8192
rect 7892 8128 7908 8192
rect 7972 8128 7988 8192
rect 8052 8128 8058 8192
rect 7742 8127 8058 8128
rect 12273 8192 12589 8193
rect 12273 8128 12279 8192
rect 12343 8128 12359 8192
rect 12423 8128 12439 8192
rect 12503 8128 12519 8192
rect 12583 8128 12589 8192
rect 12273 8127 12589 8128
rect 16804 8192 17120 8193
rect 16804 8128 16810 8192
rect 16874 8128 16890 8192
rect 16954 8128 16970 8192
rect 17034 8128 17050 8192
rect 17114 8128 17120 8192
rect 16804 8127 17120 8128
rect 3871 7648 4187 7649
rect 3871 7584 3877 7648
rect 3941 7584 3957 7648
rect 4021 7584 4037 7648
rect 4101 7584 4117 7648
rect 4181 7584 4187 7648
rect 3871 7583 4187 7584
rect 8402 7648 8718 7649
rect 8402 7584 8408 7648
rect 8472 7584 8488 7648
rect 8552 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8718 7648
rect 8402 7583 8718 7584
rect 12933 7648 13249 7649
rect 12933 7584 12939 7648
rect 13003 7584 13019 7648
rect 13083 7584 13099 7648
rect 13163 7584 13179 7648
rect 13243 7584 13249 7648
rect 12933 7583 13249 7584
rect 17464 7648 17780 7649
rect 17464 7584 17470 7648
rect 17534 7584 17550 7648
rect 17614 7584 17630 7648
rect 17694 7584 17710 7648
rect 17774 7584 17780 7648
rect 17464 7583 17780 7584
rect 3211 7104 3527 7105
rect 3211 7040 3217 7104
rect 3281 7040 3297 7104
rect 3361 7040 3377 7104
rect 3441 7040 3457 7104
rect 3521 7040 3527 7104
rect 3211 7039 3527 7040
rect 7742 7104 8058 7105
rect 7742 7040 7748 7104
rect 7812 7040 7828 7104
rect 7892 7040 7908 7104
rect 7972 7040 7988 7104
rect 8052 7040 8058 7104
rect 7742 7039 8058 7040
rect 12273 7104 12589 7105
rect 12273 7040 12279 7104
rect 12343 7040 12359 7104
rect 12423 7040 12439 7104
rect 12503 7040 12519 7104
rect 12583 7040 12589 7104
rect 12273 7039 12589 7040
rect 16804 7104 17120 7105
rect 16804 7040 16810 7104
rect 16874 7040 16890 7104
rect 16954 7040 16970 7104
rect 17034 7040 17050 7104
rect 17114 7040 17120 7104
rect 16804 7039 17120 7040
rect 3871 6560 4187 6561
rect 3871 6496 3877 6560
rect 3941 6496 3957 6560
rect 4021 6496 4037 6560
rect 4101 6496 4117 6560
rect 4181 6496 4187 6560
rect 3871 6495 4187 6496
rect 8402 6560 8718 6561
rect 8402 6496 8408 6560
rect 8472 6496 8488 6560
rect 8552 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8718 6560
rect 8402 6495 8718 6496
rect 12933 6560 13249 6561
rect 12933 6496 12939 6560
rect 13003 6496 13019 6560
rect 13083 6496 13099 6560
rect 13163 6496 13179 6560
rect 13243 6496 13249 6560
rect 12933 6495 13249 6496
rect 17464 6560 17780 6561
rect 17464 6496 17470 6560
rect 17534 6496 17550 6560
rect 17614 6496 17630 6560
rect 17694 6496 17710 6560
rect 17774 6496 17780 6560
rect 17464 6495 17780 6496
rect 3211 6016 3527 6017
rect 3211 5952 3217 6016
rect 3281 5952 3297 6016
rect 3361 5952 3377 6016
rect 3441 5952 3457 6016
rect 3521 5952 3527 6016
rect 3211 5951 3527 5952
rect 7742 6016 8058 6017
rect 7742 5952 7748 6016
rect 7812 5952 7828 6016
rect 7892 5952 7908 6016
rect 7972 5952 7988 6016
rect 8052 5952 8058 6016
rect 7742 5951 8058 5952
rect 12273 6016 12589 6017
rect 12273 5952 12279 6016
rect 12343 5952 12359 6016
rect 12423 5952 12439 6016
rect 12503 5952 12519 6016
rect 12583 5952 12589 6016
rect 12273 5951 12589 5952
rect 16804 6016 17120 6017
rect 16804 5952 16810 6016
rect 16874 5952 16890 6016
rect 16954 5952 16970 6016
rect 17034 5952 17050 6016
rect 17114 5952 17120 6016
rect 16804 5951 17120 5952
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 3871 5472 4187 5473
rect 3871 5408 3877 5472
rect 3941 5408 3957 5472
rect 4021 5408 4037 5472
rect 4101 5408 4117 5472
rect 4181 5408 4187 5472
rect 3871 5407 4187 5408
rect 8402 5472 8718 5473
rect 8402 5408 8408 5472
rect 8472 5408 8488 5472
rect 8552 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8718 5472
rect 8402 5407 8718 5408
rect 12933 5472 13249 5473
rect 12933 5408 12939 5472
rect 13003 5408 13019 5472
rect 13083 5408 13099 5472
rect 13163 5408 13179 5472
rect 13243 5408 13249 5472
rect 12933 5407 13249 5408
rect 17464 5472 17780 5473
rect 17464 5408 17470 5472
rect 17534 5408 17550 5472
rect 17614 5408 17630 5472
rect 17694 5408 17710 5472
rect 17774 5408 17780 5472
rect 17464 5407 17780 5408
rect 3211 4928 3527 4929
rect 3211 4864 3217 4928
rect 3281 4864 3297 4928
rect 3361 4864 3377 4928
rect 3441 4864 3457 4928
rect 3521 4864 3527 4928
rect 3211 4863 3527 4864
rect 7742 4928 8058 4929
rect 7742 4864 7748 4928
rect 7812 4864 7828 4928
rect 7892 4864 7908 4928
rect 7972 4864 7988 4928
rect 8052 4864 8058 4928
rect 7742 4863 8058 4864
rect 12273 4928 12589 4929
rect 12273 4864 12279 4928
rect 12343 4864 12359 4928
rect 12423 4864 12439 4928
rect 12503 4864 12519 4928
rect 12583 4864 12589 4928
rect 12273 4863 12589 4864
rect 16804 4928 17120 4929
rect 16804 4864 16810 4928
rect 16874 4864 16890 4928
rect 16954 4864 16970 4928
rect 17034 4864 17050 4928
rect 17114 4864 17120 4928
rect 16804 4863 17120 4864
rect 3871 4384 4187 4385
rect 3871 4320 3877 4384
rect 3941 4320 3957 4384
rect 4021 4320 4037 4384
rect 4101 4320 4117 4384
rect 4181 4320 4187 4384
rect 3871 4319 4187 4320
rect 8402 4384 8718 4385
rect 8402 4320 8408 4384
rect 8472 4320 8488 4384
rect 8552 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8718 4384
rect 8402 4319 8718 4320
rect 12933 4384 13249 4385
rect 12933 4320 12939 4384
rect 13003 4320 13019 4384
rect 13083 4320 13099 4384
rect 13163 4320 13179 4384
rect 13243 4320 13249 4384
rect 12933 4319 13249 4320
rect 17464 4384 17780 4385
rect 17464 4320 17470 4384
rect 17534 4320 17550 4384
rect 17614 4320 17630 4384
rect 17694 4320 17710 4384
rect 17774 4320 17780 4384
rect 17464 4319 17780 4320
rect 3211 3840 3527 3841
rect 3211 3776 3217 3840
rect 3281 3776 3297 3840
rect 3361 3776 3377 3840
rect 3441 3776 3457 3840
rect 3521 3776 3527 3840
rect 3211 3775 3527 3776
rect 7742 3840 8058 3841
rect 7742 3776 7748 3840
rect 7812 3776 7828 3840
rect 7892 3776 7908 3840
rect 7972 3776 7988 3840
rect 8052 3776 8058 3840
rect 7742 3775 8058 3776
rect 12273 3840 12589 3841
rect 12273 3776 12279 3840
rect 12343 3776 12359 3840
rect 12423 3776 12439 3840
rect 12503 3776 12519 3840
rect 12583 3776 12589 3840
rect 12273 3775 12589 3776
rect 16804 3840 17120 3841
rect 16804 3776 16810 3840
rect 16874 3776 16890 3840
rect 16954 3776 16970 3840
rect 17034 3776 17050 3840
rect 17114 3776 17120 3840
rect 16804 3775 17120 3776
rect 3871 3296 4187 3297
rect 3871 3232 3877 3296
rect 3941 3232 3957 3296
rect 4021 3232 4037 3296
rect 4101 3232 4117 3296
rect 4181 3232 4187 3296
rect 3871 3231 4187 3232
rect 8402 3296 8718 3297
rect 8402 3232 8408 3296
rect 8472 3232 8488 3296
rect 8552 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8718 3296
rect 8402 3231 8718 3232
rect 12933 3296 13249 3297
rect 12933 3232 12939 3296
rect 13003 3232 13019 3296
rect 13083 3232 13099 3296
rect 13163 3232 13179 3296
rect 13243 3232 13249 3296
rect 12933 3231 13249 3232
rect 17464 3296 17780 3297
rect 17464 3232 17470 3296
rect 17534 3232 17550 3296
rect 17614 3232 17630 3296
rect 17694 3232 17710 3296
rect 17774 3232 17780 3296
rect 17464 3231 17780 3232
rect 3211 2752 3527 2753
rect 3211 2688 3217 2752
rect 3281 2688 3297 2752
rect 3361 2688 3377 2752
rect 3441 2688 3457 2752
rect 3521 2688 3527 2752
rect 3211 2687 3527 2688
rect 7742 2752 8058 2753
rect 7742 2688 7748 2752
rect 7812 2688 7828 2752
rect 7892 2688 7908 2752
rect 7972 2688 7988 2752
rect 8052 2688 8058 2752
rect 7742 2687 8058 2688
rect 12273 2752 12589 2753
rect 12273 2688 12279 2752
rect 12343 2688 12359 2752
rect 12423 2688 12439 2752
rect 12503 2688 12519 2752
rect 12583 2688 12589 2752
rect 12273 2687 12589 2688
rect 16804 2752 17120 2753
rect 16804 2688 16810 2752
rect 16874 2688 16890 2752
rect 16954 2688 16970 2752
rect 17034 2688 17050 2752
rect 17114 2688 17120 2752
rect 16804 2687 17120 2688
rect 3871 2208 4187 2209
rect 3871 2144 3877 2208
rect 3941 2144 3957 2208
rect 4021 2144 4037 2208
rect 4101 2144 4117 2208
rect 4181 2144 4187 2208
rect 3871 2143 4187 2144
rect 8402 2208 8718 2209
rect 8402 2144 8408 2208
rect 8472 2144 8488 2208
rect 8552 2144 8568 2208
rect 8632 2144 8648 2208
rect 8712 2144 8718 2208
rect 8402 2143 8718 2144
rect 12933 2208 13249 2209
rect 12933 2144 12939 2208
rect 13003 2144 13019 2208
rect 13083 2144 13099 2208
rect 13163 2144 13179 2208
rect 13243 2144 13249 2208
rect 12933 2143 13249 2144
rect 17464 2208 17780 2209
rect 17464 2144 17470 2208
rect 17534 2144 17550 2208
rect 17614 2144 17630 2208
rect 17694 2144 17710 2208
rect 17774 2144 17780 2208
rect 17464 2143 17780 2144
<< via3 >>
rect 3217 20156 3281 20160
rect 3217 20100 3221 20156
rect 3221 20100 3277 20156
rect 3277 20100 3281 20156
rect 3217 20096 3281 20100
rect 3297 20156 3361 20160
rect 3297 20100 3301 20156
rect 3301 20100 3357 20156
rect 3357 20100 3361 20156
rect 3297 20096 3361 20100
rect 3377 20156 3441 20160
rect 3377 20100 3381 20156
rect 3381 20100 3437 20156
rect 3437 20100 3441 20156
rect 3377 20096 3441 20100
rect 3457 20156 3521 20160
rect 3457 20100 3461 20156
rect 3461 20100 3517 20156
rect 3517 20100 3521 20156
rect 3457 20096 3521 20100
rect 7748 20156 7812 20160
rect 7748 20100 7752 20156
rect 7752 20100 7808 20156
rect 7808 20100 7812 20156
rect 7748 20096 7812 20100
rect 7828 20156 7892 20160
rect 7828 20100 7832 20156
rect 7832 20100 7888 20156
rect 7888 20100 7892 20156
rect 7828 20096 7892 20100
rect 7908 20156 7972 20160
rect 7908 20100 7912 20156
rect 7912 20100 7968 20156
rect 7968 20100 7972 20156
rect 7908 20096 7972 20100
rect 7988 20156 8052 20160
rect 7988 20100 7992 20156
rect 7992 20100 8048 20156
rect 8048 20100 8052 20156
rect 7988 20096 8052 20100
rect 12279 20156 12343 20160
rect 12279 20100 12283 20156
rect 12283 20100 12339 20156
rect 12339 20100 12343 20156
rect 12279 20096 12343 20100
rect 12359 20156 12423 20160
rect 12359 20100 12363 20156
rect 12363 20100 12419 20156
rect 12419 20100 12423 20156
rect 12359 20096 12423 20100
rect 12439 20156 12503 20160
rect 12439 20100 12443 20156
rect 12443 20100 12499 20156
rect 12499 20100 12503 20156
rect 12439 20096 12503 20100
rect 12519 20156 12583 20160
rect 12519 20100 12523 20156
rect 12523 20100 12579 20156
rect 12579 20100 12583 20156
rect 12519 20096 12583 20100
rect 16810 20156 16874 20160
rect 16810 20100 16814 20156
rect 16814 20100 16870 20156
rect 16870 20100 16874 20156
rect 16810 20096 16874 20100
rect 16890 20156 16954 20160
rect 16890 20100 16894 20156
rect 16894 20100 16950 20156
rect 16950 20100 16954 20156
rect 16890 20096 16954 20100
rect 16970 20156 17034 20160
rect 16970 20100 16974 20156
rect 16974 20100 17030 20156
rect 17030 20100 17034 20156
rect 16970 20096 17034 20100
rect 17050 20156 17114 20160
rect 17050 20100 17054 20156
rect 17054 20100 17110 20156
rect 17110 20100 17114 20156
rect 17050 20096 17114 20100
rect 3877 19612 3941 19616
rect 3877 19556 3881 19612
rect 3881 19556 3937 19612
rect 3937 19556 3941 19612
rect 3877 19552 3941 19556
rect 3957 19612 4021 19616
rect 3957 19556 3961 19612
rect 3961 19556 4017 19612
rect 4017 19556 4021 19612
rect 3957 19552 4021 19556
rect 4037 19612 4101 19616
rect 4037 19556 4041 19612
rect 4041 19556 4097 19612
rect 4097 19556 4101 19612
rect 4037 19552 4101 19556
rect 4117 19612 4181 19616
rect 4117 19556 4121 19612
rect 4121 19556 4177 19612
rect 4177 19556 4181 19612
rect 4117 19552 4181 19556
rect 8408 19612 8472 19616
rect 8408 19556 8412 19612
rect 8412 19556 8468 19612
rect 8468 19556 8472 19612
rect 8408 19552 8472 19556
rect 8488 19612 8552 19616
rect 8488 19556 8492 19612
rect 8492 19556 8548 19612
rect 8548 19556 8552 19612
rect 8488 19552 8552 19556
rect 8568 19612 8632 19616
rect 8568 19556 8572 19612
rect 8572 19556 8628 19612
rect 8628 19556 8632 19612
rect 8568 19552 8632 19556
rect 8648 19612 8712 19616
rect 8648 19556 8652 19612
rect 8652 19556 8708 19612
rect 8708 19556 8712 19612
rect 8648 19552 8712 19556
rect 12939 19612 13003 19616
rect 12939 19556 12943 19612
rect 12943 19556 12999 19612
rect 12999 19556 13003 19612
rect 12939 19552 13003 19556
rect 13019 19612 13083 19616
rect 13019 19556 13023 19612
rect 13023 19556 13079 19612
rect 13079 19556 13083 19612
rect 13019 19552 13083 19556
rect 13099 19612 13163 19616
rect 13099 19556 13103 19612
rect 13103 19556 13159 19612
rect 13159 19556 13163 19612
rect 13099 19552 13163 19556
rect 13179 19612 13243 19616
rect 13179 19556 13183 19612
rect 13183 19556 13239 19612
rect 13239 19556 13243 19612
rect 13179 19552 13243 19556
rect 17470 19612 17534 19616
rect 17470 19556 17474 19612
rect 17474 19556 17530 19612
rect 17530 19556 17534 19612
rect 17470 19552 17534 19556
rect 17550 19612 17614 19616
rect 17550 19556 17554 19612
rect 17554 19556 17610 19612
rect 17610 19556 17614 19612
rect 17550 19552 17614 19556
rect 17630 19612 17694 19616
rect 17630 19556 17634 19612
rect 17634 19556 17690 19612
rect 17690 19556 17694 19612
rect 17630 19552 17694 19556
rect 17710 19612 17774 19616
rect 17710 19556 17714 19612
rect 17714 19556 17770 19612
rect 17770 19556 17774 19612
rect 17710 19552 17774 19556
rect 3217 19068 3281 19072
rect 3217 19012 3221 19068
rect 3221 19012 3277 19068
rect 3277 19012 3281 19068
rect 3217 19008 3281 19012
rect 3297 19068 3361 19072
rect 3297 19012 3301 19068
rect 3301 19012 3357 19068
rect 3357 19012 3361 19068
rect 3297 19008 3361 19012
rect 3377 19068 3441 19072
rect 3377 19012 3381 19068
rect 3381 19012 3437 19068
rect 3437 19012 3441 19068
rect 3377 19008 3441 19012
rect 3457 19068 3521 19072
rect 3457 19012 3461 19068
rect 3461 19012 3517 19068
rect 3517 19012 3521 19068
rect 3457 19008 3521 19012
rect 7748 19068 7812 19072
rect 7748 19012 7752 19068
rect 7752 19012 7808 19068
rect 7808 19012 7812 19068
rect 7748 19008 7812 19012
rect 7828 19068 7892 19072
rect 7828 19012 7832 19068
rect 7832 19012 7888 19068
rect 7888 19012 7892 19068
rect 7828 19008 7892 19012
rect 7908 19068 7972 19072
rect 7908 19012 7912 19068
rect 7912 19012 7968 19068
rect 7968 19012 7972 19068
rect 7908 19008 7972 19012
rect 7988 19068 8052 19072
rect 7988 19012 7992 19068
rect 7992 19012 8048 19068
rect 8048 19012 8052 19068
rect 7988 19008 8052 19012
rect 12279 19068 12343 19072
rect 12279 19012 12283 19068
rect 12283 19012 12339 19068
rect 12339 19012 12343 19068
rect 12279 19008 12343 19012
rect 12359 19068 12423 19072
rect 12359 19012 12363 19068
rect 12363 19012 12419 19068
rect 12419 19012 12423 19068
rect 12359 19008 12423 19012
rect 12439 19068 12503 19072
rect 12439 19012 12443 19068
rect 12443 19012 12499 19068
rect 12499 19012 12503 19068
rect 12439 19008 12503 19012
rect 12519 19068 12583 19072
rect 12519 19012 12523 19068
rect 12523 19012 12579 19068
rect 12579 19012 12583 19068
rect 12519 19008 12583 19012
rect 16810 19068 16874 19072
rect 16810 19012 16814 19068
rect 16814 19012 16870 19068
rect 16870 19012 16874 19068
rect 16810 19008 16874 19012
rect 16890 19068 16954 19072
rect 16890 19012 16894 19068
rect 16894 19012 16950 19068
rect 16950 19012 16954 19068
rect 16890 19008 16954 19012
rect 16970 19068 17034 19072
rect 16970 19012 16974 19068
rect 16974 19012 17030 19068
rect 17030 19012 17034 19068
rect 16970 19008 17034 19012
rect 17050 19068 17114 19072
rect 17050 19012 17054 19068
rect 17054 19012 17110 19068
rect 17110 19012 17114 19068
rect 17050 19008 17114 19012
rect 3877 18524 3941 18528
rect 3877 18468 3881 18524
rect 3881 18468 3937 18524
rect 3937 18468 3941 18524
rect 3877 18464 3941 18468
rect 3957 18524 4021 18528
rect 3957 18468 3961 18524
rect 3961 18468 4017 18524
rect 4017 18468 4021 18524
rect 3957 18464 4021 18468
rect 4037 18524 4101 18528
rect 4037 18468 4041 18524
rect 4041 18468 4097 18524
rect 4097 18468 4101 18524
rect 4037 18464 4101 18468
rect 4117 18524 4181 18528
rect 4117 18468 4121 18524
rect 4121 18468 4177 18524
rect 4177 18468 4181 18524
rect 4117 18464 4181 18468
rect 8408 18524 8472 18528
rect 8408 18468 8412 18524
rect 8412 18468 8468 18524
rect 8468 18468 8472 18524
rect 8408 18464 8472 18468
rect 8488 18524 8552 18528
rect 8488 18468 8492 18524
rect 8492 18468 8548 18524
rect 8548 18468 8552 18524
rect 8488 18464 8552 18468
rect 8568 18524 8632 18528
rect 8568 18468 8572 18524
rect 8572 18468 8628 18524
rect 8628 18468 8632 18524
rect 8568 18464 8632 18468
rect 8648 18524 8712 18528
rect 8648 18468 8652 18524
rect 8652 18468 8708 18524
rect 8708 18468 8712 18524
rect 8648 18464 8712 18468
rect 12939 18524 13003 18528
rect 12939 18468 12943 18524
rect 12943 18468 12999 18524
rect 12999 18468 13003 18524
rect 12939 18464 13003 18468
rect 13019 18524 13083 18528
rect 13019 18468 13023 18524
rect 13023 18468 13079 18524
rect 13079 18468 13083 18524
rect 13019 18464 13083 18468
rect 13099 18524 13163 18528
rect 13099 18468 13103 18524
rect 13103 18468 13159 18524
rect 13159 18468 13163 18524
rect 13099 18464 13163 18468
rect 13179 18524 13243 18528
rect 13179 18468 13183 18524
rect 13183 18468 13239 18524
rect 13239 18468 13243 18524
rect 13179 18464 13243 18468
rect 17470 18524 17534 18528
rect 17470 18468 17474 18524
rect 17474 18468 17530 18524
rect 17530 18468 17534 18524
rect 17470 18464 17534 18468
rect 17550 18524 17614 18528
rect 17550 18468 17554 18524
rect 17554 18468 17610 18524
rect 17610 18468 17614 18524
rect 17550 18464 17614 18468
rect 17630 18524 17694 18528
rect 17630 18468 17634 18524
rect 17634 18468 17690 18524
rect 17690 18468 17694 18524
rect 17630 18464 17694 18468
rect 17710 18524 17774 18528
rect 17710 18468 17714 18524
rect 17714 18468 17770 18524
rect 17770 18468 17774 18524
rect 17710 18464 17774 18468
rect 3217 17980 3281 17984
rect 3217 17924 3221 17980
rect 3221 17924 3277 17980
rect 3277 17924 3281 17980
rect 3217 17920 3281 17924
rect 3297 17980 3361 17984
rect 3297 17924 3301 17980
rect 3301 17924 3357 17980
rect 3357 17924 3361 17980
rect 3297 17920 3361 17924
rect 3377 17980 3441 17984
rect 3377 17924 3381 17980
rect 3381 17924 3437 17980
rect 3437 17924 3441 17980
rect 3377 17920 3441 17924
rect 3457 17980 3521 17984
rect 3457 17924 3461 17980
rect 3461 17924 3517 17980
rect 3517 17924 3521 17980
rect 3457 17920 3521 17924
rect 7748 17980 7812 17984
rect 7748 17924 7752 17980
rect 7752 17924 7808 17980
rect 7808 17924 7812 17980
rect 7748 17920 7812 17924
rect 7828 17980 7892 17984
rect 7828 17924 7832 17980
rect 7832 17924 7888 17980
rect 7888 17924 7892 17980
rect 7828 17920 7892 17924
rect 7908 17980 7972 17984
rect 7908 17924 7912 17980
rect 7912 17924 7968 17980
rect 7968 17924 7972 17980
rect 7908 17920 7972 17924
rect 7988 17980 8052 17984
rect 7988 17924 7992 17980
rect 7992 17924 8048 17980
rect 8048 17924 8052 17980
rect 7988 17920 8052 17924
rect 12279 17980 12343 17984
rect 12279 17924 12283 17980
rect 12283 17924 12339 17980
rect 12339 17924 12343 17980
rect 12279 17920 12343 17924
rect 12359 17980 12423 17984
rect 12359 17924 12363 17980
rect 12363 17924 12419 17980
rect 12419 17924 12423 17980
rect 12359 17920 12423 17924
rect 12439 17980 12503 17984
rect 12439 17924 12443 17980
rect 12443 17924 12499 17980
rect 12499 17924 12503 17980
rect 12439 17920 12503 17924
rect 12519 17980 12583 17984
rect 12519 17924 12523 17980
rect 12523 17924 12579 17980
rect 12579 17924 12583 17980
rect 12519 17920 12583 17924
rect 16810 17980 16874 17984
rect 16810 17924 16814 17980
rect 16814 17924 16870 17980
rect 16870 17924 16874 17980
rect 16810 17920 16874 17924
rect 16890 17980 16954 17984
rect 16890 17924 16894 17980
rect 16894 17924 16950 17980
rect 16950 17924 16954 17980
rect 16890 17920 16954 17924
rect 16970 17980 17034 17984
rect 16970 17924 16974 17980
rect 16974 17924 17030 17980
rect 17030 17924 17034 17980
rect 16970 17920 17034 17924
rect 17050 17980 17114 17984
rect 17050 17924 17054 17980
rect 17054 17924 17110 17980
rect 17110 17924 17114 17980
rect 17050 17920 17114 17924
rect 3877 17436 3941 17440
rect 3877 17380 3881 17436
rect 3881 17380 3937 17436
rect 3937 17380 3941 17436
rect 3877 17376 3941 17380
rect 3957 17436 4021 17440
rect 3957 17380 3961 17436
rect 3961 17380 4017 17436
rect 4017 17380 4021 17436
rect 3957 17376 4021 17380
rect 4037 17436 4101 17440
rect 4037 17380 4041 17436
rect 4041 17380 4097 17436
rect 4097 17380 4101 17436
rect 4037 17376 4101 17380
rect 4117 17436 4181 17440
rect 4117 17380 4121 17436
rect 4121 17380 4177 17436
rect 4177 17380 4181 17436
rect 4117 17376 4181 17380
rect 8408 17436 8472 17440
rect 8408 17380 8412 17436
rect 8412 17380 8468 17436
rect 8468 17380 8472 17436
rect 8408 17376 8472 17380
rect 8488 17436 8552 17440
rect 8488 17380 8492 17436
rect 8492 17380 8548 17436
rect 8548 17380 8552 17436
rect 8488 17376 8552 17380
rect 8568 17436 8632 17440
rect 8568 17380 8572 17436
rect 8572 17380 8628 17436
rect 8628 17380 8632 17436
rect 8568 17376 8632 17380
rect 8648 17436 8712 17440
rect 8648 17380 8652 17436
rect 8652 17380 8708 17436
rect 8708 17380 8712 17436
rect 8648 17376 8712 17380
rect 12939 17436 13003 17440
rect 12939 17380 12943 17436
rect 12943 17380 12999 17436
rect 12999 17380 13003 17436
rect 12939 17376 13003 17380
rect 13019 17436 13083 17440
rect 13019 17380 13023 17436
rect 13023 17380 13079 17436
rect 13079 17380 13083 17436
rect 13019 17376 13083 17380
rect 13099 17436 13163 17440
rect 13099 17380 13103 17436
rect 13103 17380 13159 17436
rect 13159 17380 13163 17436
rect 13099 17376 13163 17380
rect 13179 17436 13243 17440
rect 13179 17380 13183 17436
rect 13183 17380 13239 17436
rect 13239 17380 13243 17436
rect 13179 17376 13243 17380
rect 17470 17436 17534 17440
rect 17470 17380 17474 17436
rect 17474 17380 17530 17436
rect 17530 17380 17534 17436
rect 17470 17376 17534 17380
rect 17550 17436 17614 17440
rect 17550 17380 17554 17436
rect 17554 17380 17610 17436
rect 17610 17380 17614 17436
rect 17550 17376 17614 17380
rect 17630 17436 17694 17440
rect 17630 17380 17634 17436
rect 17634 17380 17690 17436
rect 17690 17380 17694 17436
rect 17630 17376 17694 17380
rect 17710 17436 17774 17440
rect 17710 17380 17714 17436
rect 17714 17380 17770 17436
rect 17770 17380 17774 17436
rect 17710 17376 17774 17380
rect 3217 16892 3281 16896
rect 3217 16836 3221 16892
rect 3221 16836 3277 16892
rect 3277 16836 3281 16892
rect 3217 16832 3281 16836
rect 3297 16892 3361 16896
rect 3297 16836 3301 16892
rect 3301 16836 3357 16892
rect 3357 16836 3361 16892
rect 3297 16832 3361 16836
rect 3377 16892 3441 16896
rect 3377 16836 3381 16892
rect 3381 16836 3437 16892
rect 3437 16836 3441 16892
rect 3377 16832 3441 16836
rect 3457 16892 3521 16896
rect 3457 16836 3461 16892
rect 3461 16836 3517 16892
rect 3517 16836 3521 16892
rect 3457 16832 3521 16836
rect 7748 16892 7812 16896
rect 7748 16836 7752 16892
rect 7752 16836 7808 16892
rect 7808 16836 7812 16892
rect 7748 16832 7812 16836
rect 7828 16892 7892 16896
rect 7828 16836 7832 16892
rect 7832 16836 7888 16892
rect 7888 16836 7892 16892
rect 7828 16832 7892 16836
rect 7908 16892 7972 16896
rect 7908 16836 7912 16892
rect 7912 16836 7968 16892
rect 7968 16836 7972 16892
rect 7908 16832 7972 16836
rect 7988 16892 8052 16896
rect 7988 16836 7992 16892
rect 7992 16836 8048 16892
rect 8048 16836 8052 16892
rect 7988 16832 8052 16836
rect 12279 16892 12343 16896
rect 12279 16836 12283 16892
rect 12283 16836 12339 16892
rect 12339 16836 12343 16892
rect 12279 16832 12343 16836
rect 12359 16892 12423 16896
rect 12359 16836 12363 16892
rect 12363 16836 12419 16892
rect 12419 16836 12423 16892
rect 12359 16832 12423 16836
rect 12439 16892 12503 16896
rect 12439 16836 12443 16892
rect 12443 16836 12499 16892
rect 12499 16836 12503 16892
rect 12439 16832 12503 16836
rect 12519 16892 12583 16896
rect 12519 16836 12523 16892
rect 12523 16836 12579 16892
rect 12579 16836 12583 16892
rect 12519 16832 12583 16836
rect 16810 16892 16874 16896
rect 16810 16836 16814 16892
rect 16814 16836 16870 16892
rect 16870 16836 16874 16892
rect 16810 16832 16874 16836
rect 16890 16892 16954 16896
rect 16890 16836 16894 16892
rect 16894 16836 16950 16892
rect 16950 16836 16954 16892
rect 16890 16832 16954 16836
rect 16970 16892 17034 16896
rect 16970 16836 16974 16892
rect 16974 16836 17030 16892
rect 17030 16836 17034 16892
rect 16970 16832 17034 16836
rect 17050 16892 17114 16896
rect 17050 16836 17054 16892
rect 17054 16836 17110 16892
rect 17110 16836 17114 16892
rect 17050 16832 17114 16836
rect 3877 16348 3941 16352
rect 3877 16292 3881 16348
rect 3881 16292 3937 16348
rect 3937 16292 3941 16348
rect 3877 16288 3941 16292
rect 3957 16348 4021 16352
rect 3957 16292 3961 16348
rect 3961 16292 4017 16348
rect 4017 16292 4021 16348
rect 3957 16288 4021 16292
rect 4037 16348 4101 16352
rect 4037 16292 4041 16348
rect 4041 16292 4097 16348
rect 4097 16292 4101 16348
rect 4037 16288 4101 16292
rect 4117 16348 4181 16352
rect 4117 16292 4121 16348
rect 4121 16292 4177 16348
rect 4177 16292 4181 16348
rect 4117 16288 4181 16292
rect 8408 16348 8472 16352
rect 8408 16292 8412 16348
rect 8412 16292 8468 16348
rect 8468 16292 8472 16348
rect 8408 16288 8472 16292
rect 8488 16348 8552 16352
rect 8488 16292 8492 16348
rect 8492 16292 8548 16348
rect 8548 16292 8552 16348
rect 8488 16288 8552 16292
rect 8568 16348 8632 16352
rect 8568 16292 8572 16348
rect 8572 16292 8628 16348
rect 8628 16292 8632 16348
rect 8568 16288 8632 16292
rect 8648 16348 8712 16352
rect 8648 16292 8652 16348
rect 8652 16292 8708 16348
rect 8708 16292 8712 16348
rect 8648 16288 8712 16292
rect 12939 16348 13003 16352
rect 12939 16292 12943 16348
rect 12943 16292 12999 16348
rect 12999 16292 13003 16348
rect 12939 16288 13003 16292
rect 13019 16348 13083 16352
rect 13019 16292 13023 16348
rect 13023 16292 13079 16348
rect 13079 16292 13083 16348
rect 13019 16288 13083 16292
rect 13099 16348 13163 16352
rect 13099 16292 13103 16348
rect 13103 16292 13159 16348
rect 13159 16292 13163 16348
rect 13099 16288 13163 16292
rect 13179 16348 13243 16352
rect 13179 16292 13183 16348
rect 13183 16292 13239 16348
rect 13239 16292 13243 16348
rect 13179 16288 13243 16292
rect 17470 16348 17534 16352
rect 17470 16292 17474 16348
rect 17474 16292 17530 16348
rect 17530 16292 17534 16348
rect 17470 16288 17534 16292
rect 17550 16348 17614 16352
rect 17550 16292 17554 16348
rect 17554 16292 17610 16348
rect 17610 16292 17614 16348
rect 17550 16288 17614 16292
rect 17630 16348 17694 16352
rect 17630 16292 17634 16348
rect 17634 16292 17690 16348
rect 17690 16292 17694 16348
rect 17630 16288 17694 16292
rect 17710 16348 17774 16352
rect 17710 16292 17714 16348
rect 17714 16292 17770 16348
rect 17770 16292 17774 16348
rect 17710 16288 17774 16292
rect 3217 15804 3281 15808
rect 3217 15748 3221 15804
rect 3221 15748 3277 15804
rect 3277 15748 3281 15804
rect 3217 15744 3281 15748
rect 3297 15804 3361 15808
rect 3297 15748 3301 15804
rect 3301 15748 3357 15804
rect 3357 15748 3361 15804
rect 3297 15744 3361 15748
rect 3377 15804 3441 15808
rect 3377 15748 3381 15804
rect 3381 15748 3437 15804
rect 3437 15748 3441 15804
rect 3377 15744 3441 15748
rect 3457 15804 3521 15808
rect 3457 15748 3461 15804
rect 3461 15748 3517 15804
rect 3517 15748 3521 15804
rect 3457 15744 3521 15748
rect 7748 15804 7812 15808
rect 7748 15748 7752 15804
rect 7752 15748 7808 15804
rect 7808 15748 7812 15804
rect 7748 15744 7812 15748
rect 7828 15804 7892 15808
rect 7828 15748 7832 15804
rect 7832 15748 7888 15804
rect 7888 15748 7892 15804
rect 7828 15744 7892 15748
rect 7908 15804 7972 15808
rect 7908 15748 7912 15804
rect 7912 15748 7968 15804
rect 7968 15748 7972 15804
rect 7908 15744 7972 15748
rect 7988 15804 8052 15808
rect 7988 15748 7992 15804
rect 7992 15748 8048 15804
rect 8048 15748 8052 15804
rect 7988 15744 8052 15748
rect 12279 15804 12343 15808
rect 12279 15748 12283 15804
rect 12283 15748 12339 15804
rect 12339 15748 12343 15804
rect 12279 15744 12343 15748
rect 12359 15804 12423 15808
rect 12359 15748 12363 15804
rect 12363 15748 12419 15804
rect 12419 15748 12423 15804
rect 12359 15744 12423 15748
rect 12439 15804 12503 15808
rect 12439 15748 12443 15804
rect 12443 15748 12499 15804
rect 12499 15748 12503 15804
rect 12439 15744 12503 15748
rect 12519 15804 12583 15808
rect 12519 15748 12523 15804
rect 12523 15748 12579 15804
rect 12579 15748 12583 15804
rect 12519 15744 12583 15748
rect 16810 15804 16874 15808
rect 16810 15748 16814 15804
rect 16814 15748 16870 15804
rect 16870 15748 16874 15804
rect 16810 15744 16874 15748
rect 16890 15804 16954 15808
rect 16890 15748 16894 15804
rect 16894 15748 16950 15804
rect 16950 15748 16954 15804
rect 16890 15744 16954 15748
rect 16970 15804 17034 15808
rect 16970 15748 16974 15804
rect 16974 15748 17030 15804
rect 17030 15748 17034 15804
rect 16970 15744 17034 15748
rect 17050 15804 17114 15808
rect 17050 15748 17054 15804
rect 17054 15748 17110 15804
rect 17110 15748 17114 15804
rect 17050 15744 17114 15748
rect 3877 15260 3941 15264
rect 3877 15204 3881 15260
rect 3881 15204 3937 15260
rect 3937 15204 3941 15260
rect 3877 15200 3941 15204
rect 3957 15260 4021 15264
rect 3957 15204 3961 15260
rect 3961 15204 4017 15260
rect 4017 15204 4021 15260
rect 3957 15200 4021 15204
rect 4037 15260 4101 15264
rect 4037 15204 4041 15260
rect 4041 15204 4097 15260
rect 4097 15204 4101 15260
rect 4037 15200 4101 15204
rect 4117 15260 4181 15264
rect 4117 15204 4121 15260
rect 4121 15204 4177 15260
rect 4177 15204 4181 15260
rect 4117 15200 4181 15204
rect 8408 15260 8472 15264
rect 8408 15204 8412 15260
rect 8412 15204 8468 15260
rect 8468 15204 8472 15260
rect 8408 15200 8472 15204
rect 8488 15260 8552 15264
rect 8488 15204 8492 15260
rect 8492 15204 8548 15260
rect 8548 15204 8552 15260
rect 8488 15200 8552 15204
rect 8568 15260 8632 15264
rect 8568 15204 8572 15260
rect 8572 15204 8628 15260
rect 8628 15204 8632 15260
rect 8568 15200 8632 15204
rect 8648 15260 8712 15264
rect 8648 15204 8652 15260
rect 8652 15204 8708 15260
rect 8708 15204 8712 15260
rect 8648 15200 8712 15204
rect 12939 15260 13003 15264
rect 12939 15204 12943 15260
rect 12943 15204 12999 15260
rect 12999 15204 13003 15260
rect 12939 15200 13003 15204
rect 13019 15260 13083 15264
rect 13019 15204 13023 15260
rect 13023 15204 13079 15260
rect 13079 15204 13083 15260
rect 13019 15200 13083 15204
rect 13099 15260 13163 15264
rect 13099 15204 13103 15260
rect 13103 15204 13159 15260
rect 13159 15204 13163 15260
rect 13099 15200 13163 15204
rect 13179 15260 13243 15264
rect 13179 15204 13183 15260
rect 13183 15204 13239 15260
rect 13239 15204 13243 15260
rect 13179 15200 13243 15204
rect 17470 15260 17534 15264
rect 17470 15204 17474 15260
rect 17474 15204 17530 15260
rect 17530 15204 17534 15260
rect 17470 15200 17534 15204
rect 17550 15260 17614 15264
rect 17550 15204 17554 15260
rect 17554 15204 17610 15260
rect 17610 15204 17614 15260
rect 17550 15200 17614 15204
rect 17630 15260 17694 15264
rect 17630 15204 17634 15260
rect 17634 15204 17690 15260
rect 17690 15204 17694 15260
rect 17630 15200 17694 15204
rect 17710 15260 17774 15264
rect 17710 15204 17714 15260
rect 17714 15204 17770 15260
rect 17770 15204 17774 15260
rect 17710 15200 17774 15204
rect 3217 14716 3281 14720
rect 3217 14660 3221 14716
rect 3221 14660 3277 14716
rect 3277 14660 3281 14716
rect 3217 14656 3281 14660
rect 3297 14716 3361 14720
rect 3297 14660 3301 14716
rect 3301 14660 3357 14716
rect 3357 14660 3361 14716
rect 3297 14656 3361 14660
rect 3377 14716 3441 14720
rect 3377 14660 3381 14716
rect 3381 14660 3437 14716
rect 3437 14660 3441 14716
rect 3377 14656 3441 14660
rect 3457 14716 3521 14720
rect 3457 14660 3461 14716
rect 3461 14660 3517 14716
rect 3517 14660 3521 14716
rect 3457 14656 3521 14660
rect 7748 14716 7812 14720
rect 7748 14660 7752 14716
rect 7752 14660 7808 14716
rect 7808 14660 7812 14716
rect 7748 14656 7812 14660
rect 7828 14716 7892 14720
rect 7828 14660 7832 14716
rect 7832 14660 7888 14716
rect 7888 14660 7892 14716
rect 7828 14656 7892 14660
rect 7908 14716 7972 14720
rect 7908 14660 7912 14716
rect 7912 14660 7968 14716
rect 7968 14660 7972 14716
rect 7908 14656 7972 14660
rect 7988 14716 8052 14720
rect 7988 14660 7992 14716
rect 7992 14660 8048 14716
rect 8048 14660 8052 14716
rect 7988 14656 8052 14660
rect 12279 14716 12343 14720
rect 12279 14660 12283 14716
rect 12283 14660 12339 14716
rect 12339 14660 12343 14716
rect 12279 14656 12343 14660
rect 12359 14716 12423 14720
rect 12359 14660 12363 14716
rect 12363 14660 12419 14716
rect 12419 14660 12423 14716
rect 12359 14656 12423 14660
rect 12439 14716 12503 14720
rect 12439 14660 12443 14716
rect 12443 14660 12499 14716
rect 12499 14660 12503 14716
rect 12439 14656 12503 14660
rect 12519 14716 12583 14720
rect 12519 14660 12523 14716
rect 12523 14660 12579 14716
rect 12579 14660 12583 14716
rect 12519 14656 12583 14660
rect 16810 14716 16874 14720
rect 16810 14660 16814 14716
rect 16814 14660 16870 14716
rect 16870 14660 16874 14716
rect 16810 14656 16874 14660
rect 16890 14716 16954 14720
rect 16890 14660 16894 14716
rect 16894 14660 16950 14716
rect 16950 14660 16954 14716
rect 16890 14656 16954 14660
rect 16970 14716 17034 14720
rect 16970 14660 16974 14716
rect 16974 14660 17030 14716
rect 17030 14660 17034 14716
rect 16970 14656 17034 14660
rect 17050 14716 17114 14720
rect 17050 14660 17054 14716
rect 17054 14660 17110 14716
rect 17110 14660 17114 14716
rect 17050 14656 17114 14660
rect 3877 14172 3941 14176
rect 3877 14116 3881 14172
rect 3881 14116 3937 14172
rect 3937 14116 3941 14172
rect 3877 14112 3941 14116
rect 3957 14172 4021 14176
rect 3957 14116 3961 14172
rect 3961 14116 4017 14172
rect 4017 14116 4021 14172
rect 3957 14112 4021 14116
rect 4037 14172 4101 14176
rect 4037 14116 4041 14172
rect 4041 14116 4097 14172
rect 4097 14116 4101 14172
rect 4037 14112 4101 14116
rect 4117 14172 4181 14176
rect 4117 14116 4121 14172
rect 4121 14116 4177 14172
rect 4177 14116 4181 14172
rect 4117 14112 4181 14116
rect 8408 14172 8472 14176
rect 8408 14116 8412 14172
rect 8412 14116 8468 14172
rect 8468 14116 8472 14172
rect 8408 14112 8472 14116
rect 8488 14172 8552 14176
rect 8488 14116 8492 14172
rect 8492 14116 8548 14172
rect 8548 14116 8552 14172
rect 8488 14112 8552 14116
rect 8568 14172 8632 14176
rect 8568 14116 8572 14172
rect 8572 14116 8628 14172
rect 8628 14116 8632 14172
rect 8568 14112 8632 14116
rect 8648 14172 8712 14176
rect 8648 14116 8652 14172
rect 8652 14116 8708 14172
rect 8708 14116 8712 14172
rect 8648 14112 8712 14116
rect 12939 14172 13003 14176
rect 12939 14116 12943 14172
rect 12943 14116 12999 14172
rect 12999 14116 13003 14172
rect 12939 14112 13003 14116
rect 13019 14172 13083 14176
rect 13019 14116 13023 14172
rect 13023 14116 13079 14172
rect 13079 14116 13083 14172
rect 13019 14112 13083 14116
rect 13099 14172 13163 14176
rect 13099 14116 13103 14172
rect 13103 14116 13159 14172
rect 13159 14116 13163 14172
rect 13099 14112 13163 14116
rect 13179 14172 13243 14176
rect 13179 14116 13183 14172
rect 13183 14116 13239 14172
rect 13239 14116 13243 14172
rect 13179 14112 13243 14116
rect 17470 14172 17534 14176
rect 17470 14116 17474 14172
rect 17474 14116 17530 14172
rect 17530 14116 17534 14172
rect 17470 14112 17534 14116
rect 17550 14172 17614 14176
rect 17550 14116 17554 14172
rect 17554 14116 17610 14172
rect 17610 14116 17614 14172
rect 17550 14112 17614 14116
rect 17630 14172 17694 14176
rect 17630 14116 17634 14172
rect 17634 14116 17690 14172
rect 17690 14116 17694 14172
rect 17630 14112 17694 14116
rect 17710 14172 17774 14176
rect 17710 14116 17714 14172
rect 17714 14116 17770 14172
rect 17770 14116 17774 14172
rect 17710 14112 17774 14116
rect 3217 13628 3281 13632
rect 3217 13572 3221 13628
rect 3221 13572 3277 13628
rect 3277 13572 3281 13628
rect 3217 13568 3281 13572
rect 3297 13628 3361 13632
rect 3297 13572 3301 13628
rect 3301 13572 3357 13628
rect 3357 13572 3361 13628
rect 3297 13568 3361 13572
rect 3377 13628 3441 13632
rect 3377 13572 3381 13628
rect 3381 13572 3437 13628
rect 3437 13572 3441 13628
rect 3377 13568 3441 13572
rect 3457 13628 3521 13632
rect 3457 13572 3461 13628
rect 3461 13572 3517 13628
rect 3517 13572 3521 13628
rect 3457 13568 3521 13572
rect 7748 13628 7812 13632
rect 7748 13572 7752 13628
rect 7752 13572 7808 13628
rect 7808 13572 7812 13628
rect 7748 13568 7812 13572
rect 7828 13628 7892 13632
rect 7828 13572 7832 13628
rect 7832 13572 7888 13628
rect 7888 13572 7892 13628
rect 7828 13568 7892 13572
rect 7908 13628 7972 13632
rect 7908 13572 7912 13628
rect 7912 13572 7968 13628
rect 7968 13572 7972 13628
rect 7908 13568 7972 13572
rect 7988 13628 8052 13632
rect 7988 13572 7992 13628
rect 7992 13572 8048 13628
rect 8048 13572 8052 13628
rect 7988 13568 8052 13572
rect 12279 13628 12343 13632
rect 12279 13572 12283 13628
rect 12283 13572 12339 13628
rect 12339 13572 12343 13628
rect 12279 13568 12343 13572
rect 12359 13628 12423 13632
rect 12359 13572 12363 13628
rect 12363 13572 12419 13628
rect 12419 13572 12423 13628
rect 12359 13568 12423 13572
rect 12439 13628 12503 13632
rect 12439 13572 12443 13628
rect 12443 13572 12499 13628
rect 12499 13572 12503 13628
rect 12439 13568 12503 13572
rect 12519 13628 12583 13632
rect 12519 13572 12523 13628
rect 12523 13572 12579 13628
rect 12579 13572 12583 13628
rect 12519 13568 12583 13572
rect 16810 13628 16874 13632
rect 16810 13572 16814 13628
rect 16814 13572 16870 13628
rect 16870 13572 16874 13628
rect 16810 13568 16874 13572
rect 16890 13628 16954 13632
rect 16890 13572 16894 13628
rect 16894 13572 16950 13628
rect 16950 13572 16954 13628
rect 16890 13568 16954 13572
rect 16970 13628 17034 13632
rect 16970 13572 16974 13628
rect 16974 13572 17030 13628
rect 17030 13572 17034 13628
rect 16970 13568 17034 13572
rect 17050 13628 17114 13632
rect 17050 13572 17054 13628
rect 17054 13572 17110 13628
rect 17110 13572 17114 13628
rect 17050 13568 17114 13572
rect 3877 13084 3941 13088
rect 3877 13028 3881 13084
rect 3881 13028 3937 13084
rect 3937 13028 3941 13084
rect 3877 13024 3941 13028
rect 3957 13084 4021 13088
rect 3957 13028 3961 13084
rect 3961 13028 4017 13084
rect 4017 13028 4021 13084
rect 3957 13024 4021 13028
rect 4037 13084 4101 13088
rect 4037 13028 4041 13084
rect 4041 13028 4097 13084
rect 4097 13028 4101 13084
rect 4037 13024 4101 13028
rect 4117 13084 4181 13088
rect 4117 13028 4121 13084
rect 4121 13028 4177 13084
rect 4177 13028 4181 13084
rect 4117 13024 4181 13028
rect 8408 13084 8472 13088
rect 8408 13028 8412 13084
rect 8412 13028 8468 13084
rect 8468 13028 8472 13084
rect 8408 13024 8472 13028
rect 8488 13084 8552 13088
rect 8488 13028 8492 13084
rect 8492 13028 8548 13084
rect 8548 13028 8552 13084
rect 8488 13024 8552 13028
rect 8568 13084 8632 13088
rect 8568 13028 8572 13084
rect 8572 13028 8628 13084
rect 8628 13028 8632 13084
rect 8568 13024 8632 13028
rect 8648 13084 8712 13088
rect 8648 13028 8652 13084
rect 8652 13028 8708 13084
rect 8708 13028 8712 13084
rect 8648 13024 8712 13028
rect 12939 13084 13003 13088
rect 12939 13028 12943 13084
rect 12943 13028 12999 13084
rect 12999 13028 13003 13084
rect 12939 13024 13003 13028
rect 13019 13084 13083 13088
rect 13019 13028 13023 13084
rect 13023 13028 13079 13084
rect 13079 13028 13083 13084
rect 13019 13024 13083 13028
rect 13099 13084 13163 13088
rect 13099 13028 13103 13084
rect 13103 13028 13159 13084
rect 13159 13028 13163 13084
rect 13099 13024 13163 13028
rect 13179 13084 13243 13088
rect 13179 13028 13183 13084
rect 13183 13028 13239 13084
rect 13239 13028 13243 13084
rect 13179 13024 13243 13028
rect 17470 13084 17534 13088
rect 17470 13028 17474 13084
rect 17474 13028 17530 13084
rect 17530 13028 17534 13084
rect 17470 13024 17534 13028
rect 17550 13084 17614 13088
rect 17550 13028 17554 13084
rect 17554 13028 17610 13084
rect 17610 13028 17614 13084
rect 17550 13024 17614 13028
rect 17630 13084 17694 13088
rect 17630 13028 17634 13084
rect 17634 13028 17690 13084
rect 17690 13028 17694 13084
rect 17630 13024 17694 13028
rect 17710 13084 17774 13088
rect 17710 13028 17714 13084
rect 17714 13028 17770 13084
rect 17770 13028 17774 13084
rect 17710 13024 17774 13028
rect 3217 12540 3281 12544
rect 3217 12484 3221 12540
rect 3221 12484 3277 12540
rect 3277 12484 3281 12540
rect 3217 12480 3281 12484
rect 3297 12540 3361 12544
rect 3297 12484 3301 12540
rect 3301 12484 3357 12540
rect 3357 12484 3361 12540
rect 3297 12480 3361 12484
rect 3377 12540 3441 12544
rect 3377 12484 3381 12540
rect 3381 12484 3437 12540
rect 3437 12484 3441 12540
rect 3377 12480 3441 12484
rect 3457 12540 3521 12544
rect 3457 12484 3461 12540
rect 3461 12484 3517 12540
rect 3517 12484 3521 12540
rect 3457 12480 3521 12484
rect 7748 12540 7812 12544
rect 7748 12484 7752 12540
rect 7752 12484 7808 12540
rect 7808 12484 7812 12540
rect 7748 12480 7812 12484
rect 7828 12540 7892 12544
rect 7828 12484 7832 12540
rect 7832 12484 7888 12540
rect 7888 12484 7892 12540
rect 7828 12480 7892 12484
rect 7908 12540 7972 12544
rect 7908 12484 7912 12540
rect 7912 12484 7968 12540
rect 7968 12484 7972 12540
rect 7908 12480 7972 12484
rect 7988 12540 8052 12544
rect 7988 12484 7992 12540
rect 7992 12484 8048 12540
rect 8048 12484 8052 12540
rect 7988 12480 8052 12484
rect 12279 12540 12343 12544
rect 12279 12484 12283 12540
rect 12283 12484 12339 12540
rect 12339 12484 12343 12540
rect 12279 12480 12343 12484
rect 12359 12540 12423 12544
rect 12359 12484 12363 12540
rect 12363 12484 12419 12540
rect 12419 12484 12423 12540
rect 12359 12480 12423 12484
rect 12439 12540 12503 12544
rect 12439 12484 12443 12540
rect 12443 12484 12499 12540
rect 12499 12484 12503 12540
rect 12439 12480 12503 12484
rect 12519 12540 12583 12544
rect 12519 12484 12523 12540
rect 12523 12484 12579 12540
rect 12579 12484 12583 12540
rect 12519 12480 12583 12484
rect 16810 12540 16874 12544
rect 16810 12484 16814 12540
rect 16814 12484 16870 12540
rect 16870 12484 16874 12540
rect 16810 12480 16874 12484
rect 16890 12540 16954 12544
rect 16890 12484 16894 12540
rect 16894 12484 16950 12540
rect 16950 12484 16954 12540
rect 16890 12480 16954 12484
rect 16970 12540 17034 12544
rect 16970 12484 16974 12540
rect 16974 12484 17030 12540
rect 17030 12484 17034 12540
rect 16970 12480 17034 12484
rect 17050 12540 17114 12544
rect 17050 12484 17054 12540
rect 17054 12484 17110 12540
rect 17110 12484 17114 12540
rect 17050 12480 17114 12484
rect 4292 12412 4356 12476
rect 3877 11996 3941 12000
rect 3877 11940 3881 11996
rect 3881 11940 3937 11996
rect 3937 11940 3941 11996
rect 3877 11936 3941 11940
rect 3957 11996 4021 12000
rect 3957 11940 3961 11996
rect 3961 11940 4017 11996
rect 4017 11940 4021 11996
rect 3957 11936 4021 11940
rect 4037 11996 4101 12000
rect 4037 11940 4041 11996
rect 4041 11940 4097 11996
rect 4097 11940 4101 11996
rect 4037 11936 4101 11940
rect 4117 11996 4181 12000
rect 4117 11940 4121 11996
rect 4121 11940 4177 11996
rect 4177 11940 4181 11996
rect 4117 11936 4181 11940
rect 8408 11996 8472 12000
rect 8408 11940 8412 11996
rect 8412 11940 8468 11996
rect 8468 11940 8472 11996
rect 8408 11936 8472 11940
rect 8488 11996 8552 12000
rect 8488 11940 8492 11996
rect 8492 11940 8548 11996
rect 8548 11940 8552 11996
rect 8488 11936 8552 11940
rect 8568 11996 8632 12000
rect 8568 11940 8572 11996
rect 8572 11940 8628 11996
rect 8628 11940 8632 11996
rect 8568 11936 8632 11940
rect 8648 11996 8712 12000
rect 8648 11940 8652 11996
rect 8652 11940 8708 11996
rect 8708 11940 8712 11996
rect 8648 11936 8712 11940
rect 12939 11996 13003 12000
rect 12939 11940 12943 11996
rect 12943 11940 12999 11996
rect 12999 11940 13003 11996
rect 12939 11936 13003 11940
rect 13019 11996 13083 12000
rect 13019 11940 13023 11996
rect 13023 11940 13079 11996
rect 13079 11940 13083 11996
rect 13019 11936 13083 11940
rect 13099 11996 13163 12000
rect 13099 11940 13103 11996
rect 13103 11940 13159 11996
rect 13159 11940 13163 11996
rect 13099 11936 13163 11940
rect 13179 11996 13243 12000
rect 13179 11940 13183 11996
rect 13183 11940 13239 11996
rect 13239 11940 13243 11996
rect 13179 11936 13243 11940
rect 17470 11996 17534 12000
rect 17470 11940 17474 11996
rect 17474 11940 17530 11996
rect 17530 11940 17534 11996
rect 17470 11936 17534 11940
rect 17550 11996 17614 12000
rect 17550 11940 17554 11996
rect 17554 11940 17610 11996
rect 17610 11940 17614 11996
rect 17550 11936 17614 11940
rect 17630 11996 17694 12000
rect 17630 11940 17634 11996
rect 17634 11940 17690 11996
rect 17690 11940 17694 11996
rect 17630 11936 17694 11940
rect 17710 11996 17774 12000
rect 17710 11940 17714 11996
rect 17714 11940 17770 11996
rect 17770 11940 17774 11996
rect 17710 11936 17774 11940
rect 3217 11452 3281 11456
rect 3217 11396 3221 11452
rect 3221 11396 3277 11452
rect 3277 11396 3281 11452
rect 3217 11392 3281 11396
rect 3297 11452 3361 11456
rect 3297 11396 3301 11452
rect 3301 11396 3357 11452
rect 3357 11396 3361 11452
rect 3297 11392 3361 11396
rect 3377 11452 3441 11456
rect 3377 11396 3381 11452
rect 3381 11396 3437 11452
rect 3437 11396 3441 11452
rect 3377 11392 3441 11396
rect 3457 11452 3521 11456
rect 3457 11396 3461 11452
rect 3461 11396 3517 11452
rect 3517 11396 3521 11452
rect 3457 11392 3521 11396
rect 7748 11452 7812 11456
rect 7748 11396 7752 11452
rect 7752 11396 7808 11452
rect 7808 11396 7812 11452
rect 7748 11392 7812 11396
rect 7828 11452 7892 11456
rect 7828 11396 7832 11452
rect 7832 11396 7888 11452
rect 7888 11396 7892 11452
rect 7828 11392 7892 11396
rect 7908 11452 7972 11456
rect 7908 11396 7912 11452
rect 7912 11396 7968 11452
rect 7968 11396 7972 11452
rect 7908 11392 7972 11396
rect 7988 11452 8052 11456
rect 7988 11396 7992 11452
rect 7992 11396 8048 11452
rect 8048 11396 8052 11452
rect 7988 11392 8052 11396
rect 12279 11452 12343 11456
rect 12279 11396 12283 11452
rect 12283 11396 12339 11452
rect 12339 11396 12343 11452
rect 12279 11392 12343 11396
rect 12359 11452 12423 11456
rect 12359 11396 12363 11452
rect 12363 11396 12419 11452
rect 12419 11396 12423 11452
rect 12359 11392 12423 11396
rect 12439 11452 12503 11456
rect 12439 11396 12443 11452
rect 12443 11396 12499 11452
rect 12499 11396 12503 11452
rect 12439 11392 12503 11396
rect 12519 11452 12583 11456
rect 12519 11396 12523 11452
rect 12523 11396 12579 11452
rect 12579 11396 12583 11452
rect 12519 11392 12583 11396
rect 16810 11452 16874 11456
rect 16810 11396 16814 11452
rect 16814 11396 16870 11452
rect 16870 11396 16874 11452
rect 16810 11392 16874 11396
rect 16890 11452 16954 11456
rect 16890 11396 16894 11452
rect 16894 11396 16950 11452
rect 16950 11396 16954 11452
rect 16890 11392 16954 11396
rect 16970 11452 17034 11456
rect 16970 11396 16974 11452
rect 16974 11396 17030 11452
rect 17030 11396 17034 11452
rect 16970 11392 17034 11396
rect 17050 11452 17114 11456
rect 17050 11396 17054 11452
rect 17054 11396 17110 11452
rect 17110 11396 17114 11452
rect 17050 11392 17114 11396
rect 3877 10908 3941 10912
rect 3877 10852 3881 10908
rect 3881 10852 3937 10908
rect 3937 10852 3941 10908
rect 3877 10848 3941 10852
rect 3957 10908 4021 10912
rect 3957 10852 3961 10908
rect 3961 10852 4017 10908
rect 4017 10852 4021 10908
rect 3957 10848 4021 10852
rect 4037 10908 4101 10912
rect 4037 10852 4041 10908
rect 4041 10852 4097 10908
rect 4097 10852 4101 10908
rect 4037 10848 4101 10852
rect 4117 10908 4181 10912
rect 4117 10852 4121 10908
rect 4121 10852 4177 10908
rect 4177 10852 4181 10908
rect 4117 10848 4181 10852
rect 8408 10908 8472 10912
rect 8408 10852 8412 10908
rect 8412 10852 8468 10908
rect 8468 10852 8472 10908
rect 8408 10848 8472 10852
rect 8488 10908 8552 10912
rect 8488 10852 8492 10908
rect 8492 10852 8548 10908
rect 8548 10852 8552 10908
rect 8488 10848 8552 10852
rect 8568 10908 8632 10912
rect 8568 10852 8572 10908
rect 8572 10852 8628 10908
rect 8628 10852 8632 10908
rect 8568 10848 8632 10852
rect 8648 10908 8712 10912
rect 8648 10852 8652 10908
rect 8652 10852 8708 10908
rect 8708 10852 8712 10908
rect 8648 10848 8712 10852
rect 12939 10908 13003 10912
rect 12939 10852 12943 10908
rect 12943 10852 12999 10908
rect 12999 10852 13003 10908
rect 12939 10848 13003 10852
rect 13019 10908 13083 10912
rect 13019 10852 13023 10908
rect 13023 10852 13079 10908
rect 13079 10852 13083 10908
rect 13019 10848 13083 10852
rect 13099 10908 13163 10912
rect 13099 10852 13103 10908
rect 13103 10852 13159 10908
rect 13159 10852 13163 10908
rect 13099 10848 13163 10852
rect 13179 10908 13243 10912
rect 13179 10852 13183 10908
rect 13183 10852 13239 10908
rect 13239 10852 13243 10908
rect 13179 10848 13243 10852
rect 17470 10908 17534 10912
rect 17470 10852 17474 10908
rect 17474 10852 17530 10908
rect 17530 10852 17534 10908
rect 17470 10848 17534 10852
rect 17550 10908 17614 10912
rect 17550 10852 17554 10908
rect 17554 10852 17610 10908
rect 17610 10852 17614 10908
rect 17550 10848 17614 10852
rect 17630 10908 17694 10912
rect 17630 10852 17634 10908
rect 17634 10852 17690 10908
rect 17690 10852 17694 10908
rect 17630 10848 17694 10852
rect 17710 10908 17774 10912
rect 17710 10852 17714 10908
rect 17714 10852 17770 10908
rect 17770 10852 17774 10908
rect 17710 10848 17774 10852
rect 3217 10364 3281 10368
rect 3217 10308 3221 10364
rect 3221 10308 3277 10364
rect 3277 10308 3281 10364
rect 3217 10304 3281 10308
rect 3297 10364 3361 10368
rect 3297 10308 3301 10364
rect 3301 10308 3357 10364
rect 3357 10308 3361 10364
rect 3297 10304 3361 10308
rect 3377 10364 3441 10368
rect 3377 10308 3381 10364
rect 3381 10308 3437 10364
rect 3437 10308 3441 10364
rect 3377 10304 3441 10308
rect 3457 10364 3521 10368
rect 3457 10308 3461 10364
rect 3461 10308 3517 10364
rect 3517 10308 3521 10364
rect 3457 10304 3521 10308
rect 7748 10364 7812 10368
rect 7748 10308 7752 10364
rect 7752 10308 7808 10364
rect 7808 10308 7812 10364
rect 7748 10304 7812 10308
rect 7828 10364 7892 10368
rect 7828 10308 7832 10364
rect 7832 10308 7888 10364
rect 7888 10308 7892 10364
rect 7828 10304 7892 10308
rect 7908 10364 7972 10368
rect 7908 10308 7912 10364
rect 7912 10308 7968 10364
rect 7968 10308 7972 10364
rect 7908 10304 7972 10308
rect 7988 10364 8052 10368
rect 7988 10308 7992 10364
rect 7992 10308 8048 10364
rect 8048 10308 8052 10364
rect 7988 10304 8052 10308
rect 12279 10364 12343 10368
rect 12279 10308 12283 10364
rect 12283 10308 12339 10364
rect 12339 10308 12343 10364
rect 12279 10304 12343 10308
rect 12359 10364 12423 10368
rect 12359 10308 12363 10364
rect 12363 10308 12419 10364
rect 12419 10308 12423 10364
rect 12359 10304 12423 10308
rect 12439 10364 12503 10368
rect 12439 10308 12443 10364
rect 12443 10308 12499 10364
rect 12499 10308 12503 10364
rect 12439 10304 12503 10308
rect 12519 10364 12583 10368
rect 12519 10308 12523 10364
rect 12523 10308 12579 10364
rect 12579 10308 12583 10364
rect 12519 10304 12583 10308
rect 16810 10364 16874 10368
rect 16810 10308 16814 10364
rect 16814 10308 16870 10364
rect 16870 10308 16874 10364
rect 16810 10304 16874 10308
rect 16890 10364 16954 10368
rect 16890 10308 16894 10364
rect 16894 10308 16950 10364
rect 16950 10308 16954 10364
rect 16890 10304 16954 10308
rect 16970 10364 17034 10368
rect 16970 10308 16974 10364
rect 16974 10308 17030 10364
rect 17030 10308 17034 10364
rect 16970 10304 17034 10308
rect 17050 10364 17114 10368
rect 17050 10308 17054 10364
rect 17054 10308 17110 10364
rect 17110 10308 17114 10364
rect 17050 10304 17114 10308
rect 3877 9820 3941 9824
rect 3877 9764 3881 9820
rect 3881 9764 3937 9820
rect 3937 9764 3941 9820
rect 3877 9760 3941 9764
rect 3957 9820 4021 9824
rect 3957 9764 3961 9820
rect 3961 9764 4017 9820
rect 4017 9764 4021 9820
rect 3957 9760 4021 9764
rect 4037 9820 4101 9824
rect 4037 9764 4041 9820
rect 4041 9764 4097 9820
rect 4097 9764 4101 9820
rect 4037 9760 4101 9764
rect 4117 9820 4181 9824
rect 4117 9764 4121 9820
rect 4121 9764 4177 9820
rect 4177 9764 4181 9820
rect 4117 9760 4181 9764
rect 8408 9820 8472 9824
rect 8408 9764 8412 9820
rect 8412 9764 8468 9820
rect 8468 9764 8472 9820
rect 8408 9760 8472 9764
rect 8488 9820 8552 9824
rect 8488 9764 8492 9820
rect 8492 9764 8548 9820
rect 8548 9764 8552 9820
rect 8488 9760 8552 9764
rect 8568 9820 8632 9824
rect 8568 9764 8572 9820
rect 8572 9764 8628 9820
rect 8628 9764 8632 9820
rect 8568 9760 8632 9764
rect 8648 9820 8712 9824
rect 8648 9764 8652 9820
rect 8652 9764 8708 9820
rect 8708 9764 8712 9820
rect 8648 9760 8712 9764
rect 12939 9820 13003 9824
rect 12939 9764 12943 9820
rect 12943 9764 12999 9820
rect 12999 9764 13003 9820
rect 12939 9760 13003 9764
rect 13019 9820 13083 9824
rect 13019 9764 13023 9820
rect 13023 9764 13079 9820
rect 13079 9764 13083 9820
rect 13019 9760 13083 9764
rect 13099 9820 13163 9824
rect 13099 9764 13103 9820
rect 13103 9764 13159 9820
rect 13159 9764 13163 9820
rect 13099 9760 13163 9764
rect 13179 9820 13243 9824
rect 13179 9764 13183 9820
rect 13183 9764 13239 9820
rect 13239 9764 13243 9820
rect 13179 9760 13243 9764
rect 17470 9820 17534 9824
rect 17470 9764 17474 9820
rect 17474 9764 17530 9820
rect 17530 9764 17534 9820
rect 17470 9760 17534 9764
rect 17550 9820 17614 9824
rect 17550 9764 17554 9820
rect 17554 9764 17610 9820
rect 17610 9764 17614 9820
rect 17550 9760 17614 9764
rect 17630 9820 17694 9824
rect 17630 9764 17634 9820
rect 17634 9764 17690 9820
rect 17690 9764 17694 9820
rect 17630 9760 17694 9764
rect 17710 9820 17774 9824
rect 17710 9764 17714 9820
rect 17714 9764 17770 9820
rect 17770 9764 17774 9820
rect 17710 9760 17774 9764
rect 3217 9276 3281 9280
rect 3217 9220 3221 9276
rect 3221 9220 3277 9276
rect 3277 9220 3281 9276
rect 3217 9216 3281 9220
rect 3297 9276 3361 9280
rect 3297 9220 3301 9276
rect 3301 9220 3357 9276
rect 3357 9220 3361 9276
rect 3297 9216 3361 9220
rect 3377 9276 3441 9280
rect 3377 9220 3381 9276
rect 3381 9220 3437 9276
rect 3437 9220 3441 9276
rect 3377 9216 3441 9220
rect 3457 9276 3521 9280
rect 3457 9220 3461 9276
rect 3461 9220 3517 9276
rect 3517 9220 3521 9276
rect 3457 9216 3521 9220
rect 7748 9276 7812 9280
rect 7748 9220 7752 9276
rect 7752 9220 7808 9276
rect 7808 9220 7812 9276
rect 7748 9216 7812 9220
rect 7828 9276 7892 9280
rect 7828 9220 7832 9276
rect 7832 9220 7888 9276
rect 7888 9220 7892 9276
rect 7828 9216 7892 9220
rect 7908 9276 7972 9280
rect 7908 9220 7912 9276
rect 7912 9220 7968 9276
rect 7968 9220 7972 9276
rect 7908 9216 7972 9220
rect 7988 9276 8052 9280
rect 7988 9220 7992 9276
rect 7992 9220 8048 9276
rect 8048 9220 8052 9276
rect 7988 9216 8052 9220
rect 12279 9276 12343 9280
rect 12279 9220 12283 9276
rect 12283 9220 12339 9276
rect 12339 9220 12343 9276
rect 12279 9216 12343 9220
rect 12359 9276 12423 9280
rect 12359 9220 12363 9276
rect 12363 9220 12419 9276
rect 12419 9220 12423 9276
rect 12359 9216 12423 9220
rect 12439 9276 12503 9280
rect 12439 9220 12443 9276
rect 12443 9220 12499 9276
rect 12499 9220 12503 9276
rect 12439 9216 12503 9220
rect 12519 9276 12583 9280
rect 12519 9220 12523 9276
rect 12523 9220 12579 9276
rect 12579 9220 12583 9276
rect 12519 9216 12583 9220
rect 16810 9276 16874 9280
rect 16810 9220 16814 9276
rect 16814 9220 16870 9276
rect 16870 9220 16874 9276
rect 16810 9216 16874 9220
rect 16890 9276 16954 9280
rect 16890 9220 16894 9276
rect 16894 9220 16950 9276
rect 16950 9220 16954 9276
rect 16890 9216 16954 9220
rect 16970 9276 17034 9280
rect 16970 9220 16974 9276
rect 16974 9220 17030 9276
rect 17030 9220 17034 9276
rect 16970 9216 17034 9220
rect 17050 9276 17114 9280
rect 17050 9220 17054 9276
rect 17054 9220 17110 9276
rect 17110 9220 17114 9276
rect 17050 9216 17114 9220
rect 3877 8732 3941 8736
rect 3877 8676 3881 8732
rect 3881 8676 3937 8732
rect 3937 8676 3941 8732
rect 3877 8672 3941 8676
rect 3957 8732 4021 8736
rect 3957 8676 3961 8732
rect 3961 8676 4017 8732
rect 4017 8676 4021 8732
rect 3957 8672 4021 8676
rect 4037 8732 4101 8736
rect 4037 8676 4041 8732
rect 4041 8676 4097 8732
rect 4097 8676 4101 8732
rect 4037 8672 4101 8676
rect 4117 8732 4181 8736
rect 4117 8676 4121 8732
rect 4121 8676 4177 8732
rect 4177 8676 4181 8732
rect 4117 8672 4181 8676
rect 8408 8732 8472 8736
rect 8408 8676 8412 8732
rect 8412 8676 8468 8732
rect 8468 8676 8472 8732
rect 8408 8672 8472 8676
rect 8488 8732 8552 8736
rect 8488 8676 8492 8732
rect 8492 8676 8548 8732
rect 8548 8676 8552 8732
rect 8488 8672 8552 8676
rect 8568 8732 8632 8736
rect 8568 8676 8572 8732
rect 8572 8676 8628 8732
rect 8628 8676 8632 8732
rect 8568 8672 8632 8676
rect 8648 8732 8712 8736
rect 8648 8676 8652 8732
rect 8652 8676 8708 8732
rect 8708 8676 8712 8732
rect 8648 8672 8712 8676
rect 12939 8732 13003 8736
rect 12939 8676 12943 8732
rect 12943 8676 12999 8732
rect 12999 8676 13003 8732
rect 12939 8672 13003 8676
rect 13019 8732 13083 8736
rect 13019 8676 13023 8732
rect 13023 8676 13079 8732
rect 13079 8676 13083 8732
rect 13019 8672 13083 8676
rect 13099 8732 13163 8736
rect 13099 8676 13103 8732
rect 13103 8676 13159 8732
rect 13159 8676 13163 8732
rect 13099 8672 13163 8676
rect 13179 8732 13243 8736
rect 13179 8676 13183 8732
rect 13183 8676 13239 8732
rect 13239 8676 13243 8732
rect 13179 8672 13243 8676
rect 17470 8732 17534 8736
rect 17470 8676 17474 8732
rect 17474 8676 17530 8732
rect 17530 8676 17534 8732
rect 17470 8672 17534 8676
rect 17550 8732 17614 8736
rect 17550 8676 17554 8732
rect 17554 8676 17610 8732
rect 17610 8676 17614 8732
rect 17550 8672 17614 8676
rect 17630 8732 17694 8736
rect 17630 8676 17634 8732
rect 17634 8676 17690 8732
rect 17690 8676 17694 8732
rect 17630 8672 17694 8676
rect 17710 8732 17774 8736
rect 17710 8676 17714 8732
rect 17714 8676 17770 8732
rect 17770 8676 17774 8732
rect 17710 8672 17774 8676
rect 4292 8196 4356 8260
rect 3217 8188 3281 8192
rect 3217 8132 3221 8188
rect 3221 8132 3277 8188
rect 3277 8132 3281 8188
rect 3217 8128 3281 8132
rect 3297 8188 3361 8192
rect 3297 8132 3301 8188
rect 3301 8132 3357 8188
rect 3357 8132 3361 8188
rect 3297 8128 3361 8132
rect 3377 8188 3441 8192
rect 3377 8132 3381 8188
rect 3381 8132 3437 8188
rect 3437 8132 3441 8188
rect 3377 8128 3441 8132
rect 3457 8188 3521 8192
rect 3457 8132 3461 8188
rect 3461 8132 3517 8188
rect 3517 8132 3521 8188
rect 3457 8128 3521 8132
rect 7748 8188 7812 8192
rect 7748 8132 7752 8188
rect 7752 8132 7808 8188
rect 7808 8132 7812 8188
rect 7748 8128 7812 8132
rect 7828 8188 7892 8192
rect 7828 8132 7832 8188
rect 7832 8132 7888 8188
rect 7888 8132 7892 8188
rect 7828 8128 7892 8132
rect 7908 8188 7972 8192
rect 7908 8132 7912 8188
rect 7912 8132 7968 8188
rect 7968 8132 7972 8188
rect 7908 8128 7972 8132
rect 7988 8188 8052 8192
rect 7988 8132 7992 8188
rect 7992 8132 8048 8188
rect 8048 8132 8052 8188
rect 7988 8128 8052 8132
rect 12279 8188 12343 8192
rect 12279 8132 12283 8188
rect 12283 8132 12339 8188
rect 12339 8132 12343 8188
rect 12279 8128 12343 8132
rect 12359 8188 12423 8192
rect 12359 8132 12363 8188
rect 12363 8132 12419 8188
rect 12419 8132 12423 8188
rect 12359 8128 12423 8132
rect 12439 8188 12503 8192
rect 12439 8132 12443 8188
rect 12443 8132 12499 8188
rect 12499 8132 12503 8188
rect 12439 8128 12503 8132
rect 12519 8188 12583 8192
rect 12519 8132 12523 8188
rect 12523 8132 12579 8188
rect 12579 8132 12583 8188
rect 12519 8128 12583 8132
rect 16810 8188 16874 8192
rect 16810 8132 16814 8188
rect 16814 8132 16870 8188
rect 16870 8132 16874 8188
rect 16810 8128 16874 8132
rect 16890 8188 16954 8192
rect 16890 8132 16894 8188
rect 16894 8132 16950 8188
rect 16950 8132 16954 8188
rect 16890 8128 16954 8132
rect 16970 8188 17034 8192
rect 16970 8132 16974 8188
rect 16974 8132 17030 8188
rect 17030 8132 17034 8188
rect 16970 8128 17034 8132
rect 17050 8188 17114 8192
rect 17050 8132 17054 8188
rect 17054 8132 17110 8188
rect 17110 8132 17114 8188
rect 17050 8128 17114 8132
rect 3877 7644 3941 7648
rect 3877 7588 3881 7644
rect 3881 7588 3937 7644
rect 3937 7588 3941 7644
rect 3877 7584 3941 7588
rect 3957 7644 4021 7648
rect 3957 7588 3961 7644
rect 3961 7588 4017 7644
rect 4017 7588 4021 7644
rect 3957 7584 4021 7588
rect 4037 7644 4101 7648
rect 4037 7588 4041 7644
rect 4041 7588 4097 7644
rect 4097 7588 4101 7644
rect 4037 7584 4101 7588
rect 4117 7644 4181 7648
rect 4117 7588 4121 7644
rect 4121 7588 4177 7644
rect 4177 7588 4181 7644
rect 4117 7584 4181 7588
rect 8408 7644 8472 7648
rect 8408 7588 8412 7644
rect 8412 7588 8468 7644
rect 8468 7588 8472 7644
rect 8408 7584 8472 7588
rect 8488 7644 8552 7648
rect 8488 7588 8492 7644
rect 8492 7588 8548 7644
rect 8548 7588 8552 7644
rect 8488 7584 8552 7588
rect 8568 7644 8632 7648
rect 8568 7588 8572 7644
rect 8572 7588 8628 7644
rect 8628 7588 8632 7644
rect 8568 7584 8632 7588
rect 8648 7644 8712 7648
rect 8648 7588 8652 7644
rect 8652 7588 8708 7644
rect 8708 7588 8712 7644
rect 8648 7584 8712 7588
rect 12939 7644 13003 7648
rect 12939 7588 12943 7644
rect 12943 7588 12999 7644
rect 12999 7588 13003 7644
rect 12939 7584 13003 7588
rect 13019 7644 13083 7648
rect 13019 7588 13023 7644
rect 13023 7588 13079 7644
rect 13079 7588 13083 7644
rect 13019 7584 13083 7588
rect 13099 7644 13163 7648
rect 13099 7588 13103 7644
rect 13103 7588 13159 7644
rect 13159 7588 13163 7644
rect 13099 7584 13163 7588
rect 13179 7644 13243 7648
rect 13179 7588 13183 7644
rect 13183 7588 13239 7644
rect 13239 7588 13243 7644
rect 13179 7584 13243 7588
rect 17470 7644 17534 7648
rect 17470 7588 17474 7644
rect 17474 7588 17530 7644
rect 17530 7588 17534 7644
rect 17470 7584 17534 7588
rect 17550 7644 17614 7648
rect 17550 7588 17554 7644
rect 17554 7588 17610 7644
rect 17610 7588 17614 7644
rect 17550 7584 17614 7588
rect 17630 7644 17694 7648
rect 17630 7588 17634 7644
rect 17634 7588 17690 7644
rect 17690 7588 17694 7644
rect 17630 7584 17694 7588
rect 17710 7644 17774 7648
rect 17710 7588 17714 7644
rect 17714 7588 17770 7644
rect 17770 7588 17774 7644
rect 17710 7584 17774 7588
rect 3217 7100 3281 7104
rect 3217 7044 3221 7100
rect 3221 7044 3277 7100
rect 3277 7044 3281 7100
rect 3217 7040 3281 7044
rect 3297 7100 3361 7104
rect 3297 7044 3301 7100
rect 3301 7044 3357 7100
rect 3357 7044 3361 7100
rect 3297 7040 3361 7044
rect 3377 7100 3441 7104
rect 3377 7044 3381 7100
rect 3381 7044 3437 7100
rect 3437 7044 3441 7100
rect 3377 7040 3441 7044
rect 3457 7100 3521 7104
rect 3457 7044 3461 7100
rect 3461 7044 3517 7100
rect 3517 7044 3521 7100
rect 3457 7040 3521 7044
rect 7748 7100 7812 7104
rect 7748 7044 7752 7100
rect 7752 7044 7808 7100
rect 7808 7044 7812 7100
rect 7748 7040 7812 7044
rect 7828 7100 7892 7104
rect 7828 7044 7832 7100
rect 7832 7044 7888 7100
rect 7888 7044 7892 7100
rect 7828 7040 7892 7044
rect 7908 7100 7972 7104
rect 7908 7044 7912 7100
rect 7912 7044 7968 7100
rect 7968 7044 7972 7100
rect 7908 7040 7972 7044
rect 7988 7100 8052 7104
rect 7988 7044 7992 7100
rect 7992 7044 8048 7100
rect 8048 7044 8052 7100
rect 7988 7040 8052 7044
rect 12279 7100 12343 7104
rect 12279 7044 12283 7100
rect 12283 7044 12339 7100
rect 12339 7044 12343 7100
rect 12279 7040 12343 7044
rect 12359 7100 12423 7104
rect 12359 7044 12363 7100
rect 12363 7044 12419 7100
rect 12419 7044 12423 7100
rect 12359 7040 12423 7044
rect 12439 7100 12503 7104
rect 12439 7044 12443 7100
rect 12443 7044 12499 7100
rect 12499 7044 12503 7100
rect 12439 7040 12503 7044
rect 12519 7100 12583 7104
rect 12519 7044 12523 7100
rect 12523 7044 12579 7100
rect 12579 7044 12583 7100
rect 12519 7040 12583 7044
rect 16810 7100 16874 7104
rect 16810 7044 16814 7100
rect 16814 7044 16870 7100
rect 16870 7044 16874 7100
rect 16810 7040 16874 7044
rect 16890 7100 16954 7104
rect 16890 7044 16894 7100
rect 16894 7044 16950 7100
rect 16950 7044 16954 7100
rect 16890 7040 16954 7044
rect 16970 7100 17034 7104
rect 16970 7044 16974 7100
rect 16974 7044 17030 7100
rect 17030 7044 17034 7100
rect 16970 7040 17034 7044
rect 17050 7100 17114 7104
rect 17050 7044 17054 7100
rect 17054 7044 17110 7100
rect 17110 7044 17114 7100
rect 17050 7040 17114 7044
rect 3877 6556 3941 6560
rect 3877 6500 3881 6556
rect 3881 6500 3937 6556
rect 3937 6500 3941 6556
rect 3877 6496 3941 6500
rect 3957 6556 4021 6560
rect 3957 6500 3961 6556
rect 3961 6500 4017 6556
rect 4017 6500 4021 6556
rect 3957 6496 4021 6500
rect 4037 6556 4101 6560
rect 4037 6500 4041 6556
rect 4041 6500 4097 6556
rect 4097 6500 4101 6556
rect 4037 6496 4101 6500
rect 4117 6556 4181 6560
rect 4117 6500 4121 6556
rect 4121 6500 4177 6556
rect 4177 6500 4181 6556
rect 4117 6496 4181 6500
rect 8408 6556 8472 6560
rect 8408 6500 8412 6556
rect 8412 6500 8468 6556
rect 8468 6500 8472 6556
rect 8408 6496 8472 6500
rect 8488 6556 8552 6560
rect 8488 6500 8492 6556
rect 8492 6500 8548 6556
rect 8548 6500 8552 6556
rect 8488 6496 8552 6500
rect 8568 6556 8632 6560
rect 8568 6500 8572 6556
rect 8572 6500 8628 6556
rect 8628 6500 8632 6556
rect 8568 6496 8632 6500
rect 8648 6556 8712 6560
rect 8648 6500 8652 6556
rect 8652 6500 8708 6556
rect 8708 6500 8712 6556
rect 8648 6496 8712 6500
rect 12939 6556 13003 6560
rect 12939 6500 12943 6556
rect 12943 6500 12999 6556
rect 12999 6500 13003 6556
rect 12939 6496 13003 6500
rect 13019 6556 13083 6560
rect 13019 6500 13023 6556
rect 13023 6500 13079 6556
rect 13079 6500 13083 6556
rect 13019 6496 13083 6500
rect 13099 6556 13163 6560
rect 13099 6500 13103 6556
rect 13103 6500 13159 6556
rect 13159 6500 13163 6556
rect 13099 6496 13163 6500
rect 13179 6556 13243 6560
rect 13179 6500 13183 6556
rect 13183 6500 13239 6556
rect 13239 6500 13243 6556
rect 13179 6496 13243 6500
rect 17470 6556 17534 6560
rect 17470 6500 17474 6556
rect 17474 6500 17530 6556
rect 17530 6500 17534 6556
rect 17470 6496 17534 6500
rect 17550 6556 17614 6560
rect 17550 6500 17554 6556
rect 17554 6500 17610 6556
rect 17610 6500 17614 6556
rect 17550 6496 17614 6500
rect 17630 6556 17694 6560
rect 17630 6500 17634 6556
rect 17634 6500 17690 6556
rect 17690 6500 17694 6556
rect 17630 6496 17694 6500
rect 17710 6556 17774 6560
rect 17710 6500 17714 6556
rect 17714 6500 17770 6556
rect 17770 6500 17774 6556
rect 17710 6496 17774 6500
rect 3217 6012 3281 6016
rect 3217 5956 3221 6012
rect 3221 5956 3277 6012
rect 3277 5956 3281 6012
rect 3217 5952 3281 5956
rect 3297 6012 3361 6016
rect 3297 5956 3301 6012
rect 3301 5956 3357 6012
rect 3357 5956 3361 6012
rect 3297 5952 3361 5956
rect 3377 6012 3441 6016
rect 3377 5956 3381 6012
rect 3381 5956 3437 6012
rect 3437 5956 3441 6012
rect 3377 5952 3441 5956
rect 3457 6012 3521 6016
rect 3457 5956 3461 6012
rect 3461 5956 3517 6012
rect 3517 5956 3521 6012
rect 3457 5952 3521 5956
rect 7748 6012 7812 6016
rect 7748 5956 7752 6012
rect 7752 5956 7808 6012
rect 7808 5956 7812 6012
rect 7748 5952 7812 5956
rect 7828 6012 7892 6016
rect 7828 5956 7832 6012
rect 7832 5956 7888 6012
rect 7888 5956 7892 6012
rect 7828 5952 7892 5956
rect 7908 6012 7972 6016
rect 7908 5956 7912 6012
rect 7912 5956 7968 6012
rect 7968 5956 7972 6012
rect 7908 5952 7972 5956
rect 7988 6012 8052 6016
rect 7988 5956 7992 6012
rect 7992 5956 8048 6012
rect 8048 5956 8052 6012
rect 7988 5952 8052 5956
rect 12279 6012 12343 6016
rect 12279 5956 12283 6012
rect 12283 5956 12339 6012
rect 12339 5956 12343 6012
rect 12279 5952 12343 5956
rect 12359 6012 12423 6016
rect 12359 5956 12363 6012
rect 12363 5956 12419 6012
rect 12419 5956 12423 6012
rect 12359 5952 12423 5956
rect 12439 6012 12503 6016
rect 12439 5956 12443 6012
rect 12443 5956 12499 6012
rect 12499 5956 12503 6012
rect 12439 5952 12503 5956
rect 12519 6012 12583 6016
rect 12519 5956 12523 6012
rect 12523 5956 12579 6012
rect 12579 5956 12583 6012
rect 12519 5952 12583 5956
rect 16810 6012 16874 6016
rect 16810 5956 16814 6012
rect 16814 5956 16870 6012
rect 16870 5956 16874 6012
rect 16810 5952 16874 5956
rect 16890 6012 16954 6016
rect 16890 5956 16894 6012
rect 16894 5956 16950 6012
rect 16950 5956 16954 6012
rect 16890 5952 16954 5956
rect 16970 6012 17034 6016
rect 16970 5956 16974 6012
rect 16974 5956 17030 6012
rect 17030 5956 17034 6012
rect 16970 5952 17034 5956
rect 17050 6012 17114 6016
rect 17050 5956 17054 6012
rect 17054 5956 17110 6012
rect 17110 5956 17114 6012
rect 17050 5952 17114 5956
rect 3877 5468 3941 5472
rect 3877 5412 3881 5468
rect 3881 5412 3937 5468
rect 3937 5412 3941 5468
rect 3877 5408 3941 5412
rect 3957 5468 4021 5472
rect 3957 5412 3961 5468
rect 3961 5412 4017 5468
rect 4017 5412 4021 5468
rect 3957 5408 4021 5412
rect 4037 5468 4101 5472
rect 4037 5412 4041 5468
rect 4041 5412 4097 5468
rect 4097 5412 4101 5468
rect 4037 5408 4101 5412
rect 4117 5468 4181 5472
rect 4117 5412 4121 5468
rect 4121 5412 4177 5468
rect 4177 5412 4181 5468
rect 4117 5408 4181 5412
rect 8408 5468 8472 5472
rect 8408 5412 8412 5468
rect 8412 5412 8468 5468
rect 8468 5412 8472 5468
rect 8408 5408 8472 5412
rect 8488 5468 8552 5472
rect 8488 5412 8492 5468
rect 8492 5412 8548 5468
rect 8548 5412 8552 5468
rect 8488 5408 8552 5412
rect 8568 5468 8632 5472
rect 8568 5412 8572 5468
rect 8572 5412 8628 5468
rect 8628 5412 8632 5468
rect 8568 5408 8632 5412
rect 8648 5468 8712 5472
rect 8648 5412 8652 5468
rect 8652 5412 8708 5468
rect 8708 5412 8712 5468
rect 8648 5408 8712 5412
rect 12939 5468 13003 5472
rect 12939 5412 12943 5468
rect 12943 5412 12999 5468
rect 12999 5412 13003 5468
rect 12939 5408 13003 5412
rect 13019 5468 13083 5472
rect 13019 5412 13023 5468
rect 13023 5412 13079 5468
rect 13079 5412 13083 5468
rect 13019 5408 13083 5412
rect 13099 5468 13163 5472
rect 13099 5412 13103 5468
rect 13103 5412 13159 5468
rect 13159 5412 13163 5468
rect 13099 5408 13163 5412
rect 13179 5468 13243 5472
rect 13179 5412 13183 5468
rect 13183 5412 13239 5468
rect 13239 5412 13243 5468
rect 13179 5408 13243 5412
rect 17470 5468 17534 5472
rect 17470 5412 17474 5468
rect 17474 5412 17530 5468
rect 17530 5412 17534 5468
rect 17470 5408 17534 5412
rect 17550 5468 17614 5472
rect 17550 5412 17554 5468
rect 17554 5412 17610 5468
rect 17610 5412 17614 5468
rect 17550 5408 17614 5412
rect 17630 5468 17694 5472
rect 17630 5412 17634 5468
rect 17634 5412 17690 5468
rect 17690 5412 17694 5468
rect 17630 5408 17694 5412
rect 17710 5468 17774 5472
rect 17710 5412 17714 5468
rect 17714 5412 17770 5468
rect 17770 5412 17774 5468
rect 17710 5408 17774 5412
rect 3217 4924 3281 4928
rect 3217 4868 3221 4924
rect 3221 4868 3277 4924
rect 3277 4868 3281 4924
rect 3217 4864 3281 4868
rect 3297 4924 3361 4928
rect 3297 4868 3301 4924
rect 3301 4868 3357 4924
rect 3357 4868 3361 4924
rect 3297 4864 3361 4868
rect 3377 4924 3441 4928
rect 3377 4868 3381 4924
rect 3381 4868 3437 4924
rect 3437 4868 3441 4924
rect 3377 4864 3441 4868
rect 3457 4924 3521 4928
rect 3457 4868 3461 4924
rect 3461 4868 3517 4924
rect 3517 4868 3521 4924
rect 3457 4864 3521 4868
rect 7748 4924 7812 4928
rect 7748 4868 7752 4924
rect 7752 4868 7808 4924
rect 7808 4868 7812 4924
rect 7748 4864 7812 4868
rect 7828 4924 7892 4928
rect 7828 4868 7832 4924
rect 7832 4868 7888 4924
rect 7888 4868 7892 4924
rect 7828 4864 7892 4868
rect 7908 4924 7972 4928
rect 7908 4868 7912 4924
rect 7912 4868 7968 4924
rect 7968 4868 7972 4924
rect 7908 4864 7972 4868
rect 7988 4924 8052 4928
rect 7988 4868 7992 4924
rect 7992 4868 8048 4924
rect 8048 4868 8052 4924
rect 7988 4864 8052 4868
rect 12279 4924 12343 4928
rect 12279 4868 12283 4924
rect 12283 4868 12339 4924
rect 12339 4868 12343 4924
rect 12279 4864 12343 4868
rect 12359 4924 12423 4928
rect 12359 4868 12363 4924
rect 12363 4868 12419 4924
rect 12419 4868 12423 4924
rect 12359 4864 12423 4868
rect 12439 4924 12503 4928
rect 12439 4868 12443 4924
rect 12443 4868 12499 4924
rect 12499 4868 12503 4924
rect 12439 4864 12503 4868
rect 12519 4924 12583 4928
rect 12519 4868 12523 4924
rect 12523 4868 12579 4924
rect 12579 4868 12583 4924
rect 12519 4864 12583 4868
rect 16810 4924 16874 4928
rect 16810 4868 16814 4924
rect 16814 4868 16870 4924
rect 16870 4868 16874 4924
rect 16810 4864 16874 4868
rect 16890 4924 16954 4928
rect 16890 4868 16894 4924
rect 16894 4868 16950 4924
rect 16950 4868 16954 4924
rect 16890 4864 16954 4868
rect 16970 4924 17034 4928
rect 16970 4868 16974 4924
rect 16974 4868 17030 4924
rect 17030 4868 17034 4924
rect 16970 4864 17034 4868
rect 17050 4924 17114 4928
rect 17050 4868 17054 4924
rect 17054 4868 17110 4924
rect 17110 4868 17114 4924
rect 17050 4864 17114 4868
rect 3877 4380 3941 4384
rect 3877 4324 3881 4380
rect 3881 4324 3937 4380
rect 3937 4324 3941 4380
rect 3877 4320 3941 4324
rect 3957 4380 4021 4384
rect 3957 4324 3961 4380
rect 3961 4324 4017 4380
rect 4017 4324 4021 4380
rect 3957 4320 4021 4324
rect 4037 4380 4101 4384
rect 4037 4324 4041 4380
rect 4041 4324 4097 4380
rect 4097 4324 4101 4380
rect 4037 4320 4101 4324
rect 4117 4380 4181 4384
rect 4117 4324 4121 4380
rect 4121 4324 4177 4380
rect 4177 4324 4181 4380
rect 4117 4320 4181 4324
rect 8408 4380 8472 4384
rect 8408 4324 8412 4380
rect 8412 4324 8468 4380
rect 8468 4324 8472 4380
rect 8408 4320 8472 4324
rect 8488 4380 8552 4384
rect 8488 4324 8492 4380
rect 8492 4324 8548 4380
rect 8548 4324 8552 4380
rect 8488 4320 8552 4324
rect 8568 4380 8632 4384
rect 8568 4324 8572 4380
rect 8572 4324 8628 4380
rect 8628 4324 8632 4380
rect 8568 4320 8632 4324
rect 8648 4380 8712 4384
rect 8648 4324 8652 4380
rect 8652 4324 8708 4380
rect 8708 4324 8712 4380
rect 8648 4320 8712 4324
rect 12939 4380 13003 4384
rect 12939 4324 12943 4380
rect 12943 4324 12999 4380
rect 12999 4324 13003 4380
rect 12939 4320 13003 4324
rect 13019 4380 13083 4384
rect 13019 4324 13023 4380
rect 13023 4324 13079 4380
rect 13079 4324 13083 4380
rect 13019 4320 13083 4324
rect 13099 4380 13163 4384
rect 13099 4324 13103 4380
rect 13103 4324 13159 4380
rect 13159 4324 13163 4380
rect 13099 4320 13163 4324
rect 13179 4380 13243 4384
rect 13179 4324 13183 4380
rect 13183 4324 13239 4380
rect 13239 4324 13243 4380
rect 13179 4320 13243 4324
rect 17470 4380 17534 4384
rect 17470 4324 17474 4380
rect 17474 4324 17530 4380
rect 17530 4324 17534 4380
rect 17470 4320 17534 4324
rect 17550 4380 17614 4384
rect 17550 4324 17554 4380
rect 17554 4324 17610 4380
rect 17610 4324 17614 4380
rect 17550 4320 17614 4324
rect 17630 4380 17694 4384
rect 17630 4324 17634 4380
rect 17634 4324 17690 4380
rect 17690 4324 17694 4380
rect 17630 4320 17694 4324
rect 17710 4380 17774 4384
rect 17710 4324 17714 4380
rect 17714 4324 17770 4380
rect 17770 4324 17774 4380
rect 17710 4320 17774 4324
rect 3217 3836 3281 3840
rect 3217 3780 3221 3836
rect 3221 3780 3277 3836
rect 3277 3780 3281 3836
rect 3217 3776 3281 3780
rect 3297 3836 3361 3840
rect 3297 3780 3301 3836
rect 3301 3780 3357 3836
rect 3357 3780 3361 3836
rect 3297 3776 3361 3780
rect 3377 3836 3441 3840
rect 3377 3780 3381 3836
rect 3381 3780 3437 3836
rect 3437 3780 3441 3836
rect 3377 3776 3441 3780
rect 3457 3836 3521 3840
rect 3457 3780 3461 3836
rect 3461 3780 3517 3836
rect 3517 3780 3521 3836
rect 3457 3776 3521 3780
rect 7748 3836 7812 3840
rect 7748 3780 7752 3836
rect 7752 3780 7808 3836
rect 7808 3780 7812 3836
rect 7748 3776 7812 3780
rect 7828 3836 7892 3840
rect 7828 3780 7832 3836
rect 7832 3780 7888 3836
rect 7888 3780 7892 3836
rect 7828 3776 7892 3780
rect 7908 3836 7972 3840
rect 7908 3780 7912 3836
rect 7912 3780 7968 3836
rect 7968 3780 7972 3836
rect 7908 3776 7972 3780
rect 7988 3836 8052 3840
rect 7988 3780 7992 3836
rect 7992 3780 8048 3836
rect 8048 3780 8052 3836
rect 7988 3776 8052 3780
rect 12279 3836 12343 3840
rect 12279 3780 12283 3836
rect 12283 3780 12339 3836
rect 12339 3780 12343 3836
rect 12279 3776 12343 3780
rect 12359 3836 12423 3840
rect 12359 3780 12363 3836
rect 12363 3780 12419 3836
rect 12419 3780 12423 3836
rect 12359 3776 12423 3780
rect 12439 3836 12503 3840
rect 12439 3780 12443 3836
rect 12443 3780 12499 3836
rect 12499 3780 12503 3836
rect 12439 3776 12503 3780
rect 12519 3836 12583 3840
rect 12519 3780 12523 3836
rect 12523 3780 12579 3836
rect 12579 3780 12583 3836
rect 12519 3776 12583 3780
rect 16810 3836 16874 3840
rect 16810 3780 16814 3836
rect 16814 3780 16870 3836
rect 16870 3780 16874 3836
rect 16810 3776 16874 3780
rect 16890 3836 16954 3840
rect 16890 3780 16894 3836
rect 16894 3780 16950 3836
rect 16950 3780 16954 3836
rect 16890 3776 16954 3780
rect 16970 3836 17034 3840
rect 16970 3780 16974 3836
rect 16974 3780 17030 3836
rect 17030 3780 17034 3836
rect 16970 3776 17034 3780
rect 17050 3836 17114 3840
rect 17050 3780 17054 3836
rect 17054 3780 17110 3836
rect 17110 3780 17114 3836
rect 17050 3776 17114 3780
rect 3877 3292 3941 3296
rect 3877 3236 3881 3292
rect 3881 3236 3937 3292
rect 3937 3236 3941 3292
rect 3877 3232 3941 3236
rect 3957 3292 4021 3296
rect 3957 3236 3961 3292
rect 3961 3236 4017 3292
rect 4017 3236 4021 3292
rect 3957 3232 4021 3236
rect 4037 3292 4101 3296
rect 4037 3236 4041 3292
rect 4041 3236 4097 3292
rect 4097 3236 4101 3292
rect 4037 3232 4101 3236
rect 4117 3292 4181 3296
rect 4117 3236 4121 3292
rect 4121 3236 4177 3292
rect 4177 3236 4181 3292
rect 4117 3232 4181 3236
rect 8408 3292 8472 3296
rect 8408 3236 8412 3292
rect 8412 3236 8468 3292
rect 8468 3236 8472 3292
rect 8408 3232 8472 3236
rect 8488 3292 8552 3296
rect 8488 3236 8492 3292
rect 8492 3236 8548 3292
rect 8548 3236 8552 3292
rect 8488 3232 8552 3236
rect 8568 3292 8632 3296
rect 8568 3236 8572 3292
rect 8572 3236 8628 3292
rect 8628 3236 8632 3292
rect 8568 3232 8632 3236
rect 8648 3292 8712 3296
rect 8648 3236 8652 3292
rect 8652 3236 8708 3292
rect 8708 3236 8712 3292
rect 8648 3232 8712 3236
rect 12939 3292 13003 3296
rect 12939 3236 12943 3292
rect 12943 3236 12999 3292
rect 12999 3236 13003 3292
rect 12939 3232 13003 3236
rect 13019 3292 13083 3296
rect 13019 3236 13023 3292
rect 13023 3236 13079 3292
rect 13079 3236 13083 3292
rect 13019 3232 13083 3236
rect 13099 3292 13163 3296
rect 13099 3236 13103 3292
rect 13103 3236 13159 3292
rect 13159 3236 13163 3292
rect 13099 3232 13163 3236
rect 13179 3292 13243 3296
rect 13179 3236 13183 3292
rect 13183 3236 13239 3292
rect 13239 3236 13243 3292
rect 13179 3232 13243 3236
rect 17470 3292 17534 3296
rect 17470 3236 17474 3292
rect 17474 3236 17530 3292
rect 17530 3236 17534 3292
rect 17470 3232 17534 3236
rect 17550 3292 17614 3296
rect 17550 3236 17554 3292
rect 17554 3236 17610 3292
rect 17610 3236 17614 3292
rect 17550 3232 17614 3236
rect 17630 3292 17694 3296
rect 17630 3236 17634 3292
rect 17634 3236 17690 3292
rect 17690 3236 17694 3292
rect 17630 3232 17694 3236
rect 17710 3292 17774 3296
rect 17710 3236 17714 3292
rect 17714 3236 17770 3292
rect 17770 3236 17774 3292
rect 17710 3232 17774 3236
rect 3217 2748 3281 2752
rect 3217 2692 3221 2748
rect 3221 2692 3277 2748
rect 3277 2692 3281 2748
rect 3217 2688 3281 2692
rect 3297 2748 3361 2752
rect 3297 2692 3301 2748
rect 3301 2692 3357 2748
rect 3357 2692 3361 2748
rect 3297 2688 3361 2692
rect 3377 2748 3441 2752
rect 3377 2692 3381 2748
rect 3381 2692 3437 2748
rect 3437 2692 3441 2748
rect 3377 2688 3441 2692
rect 3457 2748 3521 2752
rect 3457 2692 3461 2748
rect 3461 2692 3517 2748
rect 3517 2692 3521 2748
rect 3457 2688 3521 2692
rect 7748 2748 7812 2752
rect 7748 2692 7752 2748
rect 7752 2692 7808 2748
rect 7808 2692 7812 2748
rect 7748 2688 7812 2692
rect 7828 2748 7892 2752
rect 7828 2692 7832 2748
rect 7832 2692 7888 2748
rect 7888 2692 7892 2748
rect 7828 2688 7892 2692
rect 7908 2748 7972 2752
rect 7908 2692 7912 2748
rect 7912 2692 7968 2748
rect 7968 2692 7972 2748
rect 7908 2688 7972 2692
rect 7988 2748 8052 2752
rect 7988 2692 7992 2748
rect 7992 2692 8048 2748
rect 8048 2692 8052 2748
rect 7988 2688 8052 2692
rect 12279 2748 12343 2752
rect 12279 2692 12283 2748
rect 12283 2692 12339 2748
rect 12339 2692 12343 2748
rect 12279 2688 12343 2692
rect 12359 2748 12423 2752
rect 12359 2692 12363 2748
rect 12363 2692 12419 2748
rect 12419 2692 12423 2748
rect 12359 2688 12423 2692
rect 12439 2748 12503 2752
rect 12439 2692 12443 2748
rect 12443 2692 12499 2748
rect 12499 2692 12503 2748
rect 12439 2688 12503 2692
rect 12519 2748 12583 2752
rect 12519 2692 12523 2748
rect 12523 2692 12579 2748
rect 12579 2692 12583 2748
rect 12519 2688 12583 2692
rect 16810 2748 16874 2752
rect 16810 2692 16814 2748
rect 16814 2692 16870 2748
rect 16870 2692 16874 2748
rect 16810 2688 16874 2692
rect 16890 2748 16954 2752
rect 16890 2692 16894 2748
rect 16894 2692 16950 2748
rect 16950 2692 16954 2748
rect 16890 2688 16954 2692
rect 16970 2748 17034 2752
rect 16970 2692 16974 2748
rect 16974 2692 17030 2748
rect 17030 2692 17034 2748
rect 16970 2688 17034 2692
rect 17050 2748 17114 2752
rect 17050 2692 17054 2748
rect 17054 2692 17110 2748
rect 17110 2692 17114 2748
rect 17050 2688 17114 2692
rect 3877 2204 3941 2208
rect 3877 2148 3881 2204
rect 3881 2148 3937 2204
rect 3937 2148 3941 2204
rect 3877 2144 3941 2148
rect 3957 2204 4021 2208
rect 3957 2148 3961 2204
rect 3961 2148 4017 2204
rect 4017 2148 4021 2204
rect 3957 2144 4021 2148
rect 4037 2204 4101 2208
rect 4037 2148 4041 2204
rect 4041 2148 4097 2204
rect 4097 2148 4101 2204
rect 4037 2144 4101 2148
rect 4117 2204 4181 2208
rect 4117 2148 4121 2204
rect 4121 2148 4177 2204
rect 4177 2148 4181 2204
rect 4117 2144 4181 2148
rect 8408 2204 8472 2208
rect 8408 2148 8412 2204
rect 8412 2148 8468 2204
rect 8468 2148 8472 2204
rect 8408 2144 8472 2148
rect 8488 2204 8552 2208
rect 8488 2148 8492 2204
rect 8492 2148 8548 2204
rect 8548 2148 8552 2204
rect 8488 2144 8552 2148
rect 8568 2204 8632 2208
rect 8568 2148 8572 2204
rect 8572 2148 8628 2204
rect 8628 2148 8632 2204
rect 8568 2144 8632 2148
rect 8648 2204 8712 2208
rect 8648 2148 8652 2204
rect 8652 2148 8708 2204
rect 8708 2148 8712 2204
rect 8648 2144 8712 2148
rect 12939 2204 13003 2208
rect 12939 2148 12943 2204
rect 12943 2148 12999 2204
rect 12999 2148 13003 2204
rect 12939 2144 13003 2148
rect 13019 2204 13083 2208
rect 13019 2148 13023 2204
rect 13023 2148 13079 2204
rect 13079 2148 13083 2204
rect 13019 2144 13083 2148
rect 13099 2204 13163 2208
rect 13099 2148 13103 2204
rect 13103 2148 13159 2204
rect 13159 2148 13163 2204
rect 13099 2144 13163 2148
rect 13179 2204 13243 2208
rect 13179 2148 13183 2204
rect 13183 2148 13239 2204
rect 13239 2148 13243 2204
rect 13179 2144 13243 2148
rect 17470 2204 17534 2208
rect 17470 2148 17474 2204
rect 17474 2148 17530 2204
rect 17530 2148 17534 2204
rect 17470 2144 17534 2148
rect 17550 2204 17614 2208
rect 17550 2148 17554 2204
rect 17554 2148 17610 2204
rect 17610 2148 17614 2204
rect 17550 2144 17614 2148
rect 17630 2204 17694 2208
rect 17630 2148 17634 2204
rect 17634 2148 17690 2204
rect 17690 2148 17694 2204
rect 17630 2144 17694 2148
rect 17710 2204 17774 2208
rect 17710 2148 17714 2204
rect 17714 2148 17770 2204
rect 17770 2148 17774 2204
rect 17710 2144 17774 2148
<< metal4 >>
rect 3209 20160 3529 20176
rect 3209 20096 3217 20160
rect 3281 20096 3297 20160
rect 3361 20096 3377 20160
rect 3441 20096 3457 20160
rect 3521 20096 3529 20160
rect 3209 19072 3529 20096
rect 3209 19008 3217 19072
rect 3281 19008 3297 19072
rect 3361 19008 3377 19072
rect 3441 19008 3457 19072
rect 3521 19008 3529 19072
rect 3209 18002 3529 19008
rect 3209 17984 3251 18002
rect 3487 17984 3529 18002
rect 3209 17920 3217 17984
rect 3521 17920 3529 17984
rect 3209 17766 3251 17920
rect 3487 17766 3529 17920
rect 3209 16896 3529 17766
rect 3209 16832 3217 16896
rect 3281 16832 3297 16896
rect 3361 16832 3377 16896
rect 3441 16832 3457 16896
rect 3521 16832 3529 16896
rect 3209 15808 3529 16832
rect 3209 15744 3217 15808
rect 3281 15744 3297 15808
rect 3361 15744 3377 15808
rect 3441 15744 3457 15808
rect 3521 15744 3529 15808
rect 3209 14720 3529 15744
rect 3209 14656 3217 14720
rect 3281 14656 3297 14720
rect 3361 14656 3377 14720
rect 3441 14656 3457 14720
rect 3521 14656 3529 14720
rect 3209 13632 3529 14656
rect 3209 13568 3217 13632
rect 3281 13568 3297 13632
rect 3361 13568 3377 13632
rect 3441 13568 3457 13632
rect 3521 13568 3529 13632
rect 3209 13514 3529 13568
rect 3209 13278 3251 13514
rect 3487 13278 3529 13514
rect 3209 12544 3529 13278
rect 3209 12480 3217 12544
rect 3281 12480 3297 12544
rect 3361 12480 3377 12544
rect 3441 12480 3457 12544
rect 3521 12480 3529 12544
rect 3209 11456 3529 12480
rect 3209 11392 3217 11456
rect 3281 11392 3297 11456
rect 3361 11392 3377 11456
rect 3441 11392 3457 11456
rect 3521 11392 3529 11456
rect 3209 10368 3529 11392
rect 3209 10304 3217 10368
rect 3281 10304 3297 10368
rect 3361 10304 3377 10368
rect 3441 10304 3457 10368
rect 3521 10304 3529 10368
rect 3209 9280 3529 10304
rect 3209 9216 3217 9280
rect 3281 9216 3297 9280
rect 3361 9216 3377 9280
rect 3441 9216 3457 9280
rect 3521 9216 3529 9280
rect 3209 9026 3529 9216
rect 3209 8790 3251 9026
rect 3487 8790 3529 9026
rect 3209 8192 3529 8790
rect 3209 8128 3217 8192
rect 3281 8128 3297 8192
rect 3361 8128 3377 8192
rect 3441 8128 3457 8192
rect 3521 8128 3529 8192
rect 3209 7104 3529 8128
rect 3209 7040 3217 7104
rect 3281 7040 3297 7104
rect 3361 7040 3377 7104
rect 3441 7040 3457 7104
rect 3521 7040 3529 7104
rect 3209 6016 3529 7040
rect 3209 5952 3217 6016
rect 3281 5952 3297 6016
rect 3361 5952 3377 6016
rect 3441 5952 3457 6016
rect 3521 5952 3529 6016
rect 3209 4928 3529 5952
rect 3209 4864 3217 4928
rect 3281 4864 3297 4928
rect 3361 4864 3377 4928
rect 3441 4864 3457 4928
rect 3521 4864 3529 4928
rect 3209 4538 3529 4864
rect 3209 4302 3251 4538
rect 3487 4302 3529 4538
rect 3209 3840 3529 4302
rect 3209 3776 3217 3840
rect 3281 3776 3297 3840
rect 3361 3776 3377 3840
rect 3441 3776 3457 3840
rect 3521 3776 3529 3840
rect 3209 2752 3529 3776
rect 3209 2688 3217 2752
rect 3281 2688 3297 2752
rect 3361 2688 3377 2752
rect 3441 2688 3457 2752
rect 3521 2688 3529 2752
rect 3209 2128 3529 2688
rect 3869 19616 4189 20176
rect 3869 19552 3877 19616
rect 3941 19552 3957 19616
rect 4021 19552 4037 19616
rect 4101 19552 4117 19616
rect 4181 19552 4189 19616
rect 3869 18662 4189 19552
rect 3869 18528 3911 18662
rect 4147 18528 4189 18662
rect 3869 18464 3877 18528
rect 4181 18464 4189 18528
rect 3869 18426 3911 18464
rect 4147 18426 4189 18464
rect 3869 17440 4189 18426
rect 3869 17376 3877 17440
rect 3941 17376 3957 17440
rect 4021 17376 4037 17440
rect 4101 17376 4117 17440
rect 4181 17376 4189 17440
rect 3869 16352 4189 17376
rect 3869 16288 3877 16352
rect 3941 16288 3957 16352
rect 4021 16288 4037 16352
rect 4101 16288 4117 16352
rect 4181 16288 4189 16352
rect 3869 15264 4189 16288
rect 3869 15200 3877 15264
rect 3941 15200 3957 15264
rect 4021 15200 4037 15264
rect 4101 15200 4117 15264
rect 4181 15200 4189 15264
rect 3869 14176 4189 15200
rect 3869 14112 3877 14176
rect 3941 14174 3957 14176
rect 4021 14174 4037 14176
rect 4101 14174 4117 14176
rect 4181 14112 4189 14176
rect 3869 13938 3911 14112
rect 4147 13938 4189 14112
rect 3869 13088 4189 13938
rect 3869 13024 3877 13088
rect 3941 13024 3957 13088
rect 4021 13024 4037 13088
rect 4101 13024 4117 13088
rect 4181 13024 4189 13088
rect 3869 12000 4189 13024
rect 7740 20160 8060 20176
rect 7740 20096 7748 20160
rect 7812 20096 7828 20160
rect 7892 20096 7908 20160
rect 7972 20096 7988 20160
rect 8052 20096 8060 20160
rect 7740 19072 8060 20096
rect 7740 19008 7748 19072
rect 7812 19008 7828 19072
rect 7892 19008 7908 19072
rect 7972 19008 7988 19072
rect 8052 19008 8060 19072
rect 7740 18002 8060 19008
rect 7740 17984 7782 18002
rect 8018 17984 8060 18002
rect 7740 17920 7748 17984
rect 8052 17920 8060 17984
rect 7740 17766 7782 17920
rect 8018 17766 8060 17920
rect 7740 16896 8060 17766
rect 7740 16832 7748 16896
rect 7812 16832 7828 16896
rect 7892 16832 7908 16896
rect 7972 16832 7988 16896
rect 8052 16832 8060 16896
rect 7740 15808 8060 16832
rect 7740 15744 7748 15808
rect 7812 15744 7828 15808
rect 7892 15744 7908 15808
rect 7972 15744 7988 15808
rect 8052 15744 8060 15808
rect 7740 14720 8060 15744
rect 7740 14656 7748 14720
rect 7812 14656 7828 14720
rect 7892 14656 7908 14720
rect 7972 14656 7988 14720
rect 8052 14656 8060 14720
rect 7740 13632 8060 14656
rect 7740 13568 7748 13632
rect 7812 13568 7828 13632
rect 7892 13568 7908 13632
rect 7972 13568 7988 13632
rect 8052 13568 8060 13632
rect 7740 13514 8060 13568
rect 7740 13278 7782 13514
rect 8018 13278 8060 13514
rect 7740 12544 8060 13278
rect 7740 12480 7748 12544
rect 7812 12480 7828 12544
rect 7892 12480 7908 12544
rect 7972 12480 7988 12544
rect 8052 12480 8060 12544
rect 4291 12476 4357 12477
rect 4291 12412 4292 12476
rect 4356 12412 4357 12476
rect 4291 12411 4357 12412
rect 3869 11936 3877 12000
rect 3941 11936 3957 12000
rect 4021 11936 4037 12000
rect 4101 11936 4117 12000
rect 4181 11936 4189 12000
rect 3869 10912 4189 11936
rect 3869 10848 3877 10912
rect 3941 10848 3957 10912
rect 4021 10848 4037 10912
rect 4101 10848 4117 10912
rect 4181 10848 4189 10912
rect 3869 9824 4189 10848
rect 3869 9760 3877 9824
rect 3941 9760 3957 9824
rect 4021 9760 4037 9824
rect 4101 9760 4117 9824
rect 4181 9760 4189 9824
rect 3869 9686 4189 9760
rect 3869 9450 3911 9686
rect 4147 9450 4189 9686
rect 3869 8736 4189 9450
rect 3869 8672 3877 8736
rect 3941 8672 3957 8736
rect 4021 8672 4037 8736
rect 4101 8672 4117 8736
rect 4181 8672 4189 8736
rect 3869 7648 4189 8672
rect 4294 8261 4354 12411
rect 7740 11456 8060 12480
rect 7740 11392 7748 11456
rect 7812 11392 7828 11456
rect 7892 11392 7908 11456
rect 7972 11392 7988 11456
rect 8052 11392 8060 11456
rect 7740 10368 8060 11392
rect 7740 10304 7748 10368
rect 7812 10304 7828 10368
rect 7892 10304 7908 10368
rect 7972 10304 7988 10368
rect 8052 10304 8060 10368
rect 7740 9280 8060 10304
rect 7740 9216 7748 9280
rect 7812 9216 7828 9280
rect 7892 9216 7908 9280
rect 7972 9216 7988 9280
rect 8052 9216 8060 9280
rect 7740 9026 8060 9216
rect 7740 8790 7782 9026
rect 8018 8790 8060 9026
rect 4291 8260 4357 8261
rect 4291 8196 4292 8260
rect 4356 8196 4357 8260
rect 4291 8195 4357 8196
rect 3869 7584 3877 7648
rect 3941 7584 3957 7648
rect 4021 7584 4037 7648
rect 4101 7584 4117 7648
rect 4181 7584 4189 7648
rect 3869 6560 4189 7584
rect 3869 6496 3877 6560
rect 3941 6496 3957 6560
rect 4021 6496 4037 6560
rect 4101 6496 4117 6560
rect 4181 6496 4189 6560
rect 3869 5472 4189 6496
rect 3869 5408 3877 5472
rect 3941 5408 3957 5472
rect 4021 5408 4037 5472
rect 4101 5408 4117 5472
rect 4181 5408 4189 5472
rect 3869 5198 4189 5408
rect 3869 4962 3911 5198
rect 4147 4962 4189 5198
rect 3869 4384 4189 4962
rect 3869 4320 3877 4384
rect 3941 4320 3957 4384
rect 4021 4320 4037 4384
rect 4101 4320 4117 4384
rect 4181 4320 4189 4384
rect 3869 3296 4189 4320
rect 3869 3232 3877 3296
rect 3941 3232 3957 3296
rect 4021 3232 4037 3296
rect 4101 3232 4117 3296
rect 4181 3232 4189 3296
rect 3869 2208 4189 3232
rect 3869 2144 3877 2208
rect 3941 2144 3957 2208
rect 4021 2144 4037 2208
rect 4101 2144 4117 2208
rect 4181 2144 4189 2208
rect 3869 2128 4189 2144
rect 7740 8192 8060 8790
rect 7740 8128 7748 8192
rect 7812 8128 7828 8192
rect 7892 8128 7908 8192
rect 7972 8128 7988 8192
rect 8052 8128 8060 8192
rect 7740 7104 8060 8128
rect 7740 7040 7748 7104
rect 7812 7040 7828 7104
rect 7892 7040 7908 7104
rect 7972 7040 7988 7104
rect 8052 7040 8060 7104
rect 7740 6016 8060 7040
rect 7740 5952 7748 6016
rect 7812 5952 7828 6016
rect 7892 5952 7908 6016
rect 7972 5952 7988 6016
rect 8052 5952 8060 6016
rect 7740 4928 8060 5952
rect 7740 4864 7748 4928
rect 7812 4864 7828 4928
rect 7892 4864 7908 4928
rect 7972 4864 7988 4928
rect 8052 4864 8060 4928
rect 7740 4538 8060 4864
rect 7740 4302 7782 4538
rect 8018 4302 8060 4538
rect 7740 3840 8060 4302
rect 7740 3776 7748 3840
rect 7812 3776 7828 3840
rect 7892 3776 7908 3840
rect 7972 3776 7988 3840
rect 8052 3776 8060 3840
rect 7740 2752 8060 3776
rect 7740 2688 7748 2752
rect 7812 2688 7828 2752
rect 7892 2688 7908 2752
rect 7972 2688 7988 2752
rect 8052 2688 8060 2752
rect 7740 2128 8060 2688
rect 8400 19616 8720 20176
rect 8400 19552 8408 19616
rect 8472 19552 8488 19616
rect 8552 19552 8568 19616
rect 8632 19552 8648 19616
rect 8712 19552 8720 19616
rect 8400 18662 8720 19552
rect 8400 18528 8442 18662
rect 8678 18528 8720 18662
rect 8400 18464 8408 18528
rect 8712 18464 8720 18528
rect 8400 18426 8442 18464
rect 8678 18426 8720 18464
rect 8400 17440 8720 18426
rect 8400 17376 8408 17440
rect 8472 17376 8488 17440
rect 8552 17376 8568 17440
rect 8632 17376 8648 17440
rect 8712 17376 8720 17440
rect 8400 16352 8720 17376
rect 8400 16288 8408 16352
rect 8472 16288 8488 16352
rect 8552 16288 8568 16352
rect 8632 16288 8648 16352
rect 8712 16288 8720 16352
rect 8400 15264 8720 16288
rect 8400 15200 8408 15264
rect 8472 15200 8488 15264
rect 8552 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8720 15264
rect 8400 14176 8720 15200
rect 8400 14112 8408 14176
rect 8472 14174 8488 14176
rect 8552 14174 8568 14176
rect 8632 14174 8648 14176
rect 8712 14112 8720 14176
rect 8400 13938 8442 14112
rect 8678 13938 8720 14112
rect 8400 13088 8720 13938
rect 8400 13024 8408 13088
rect 8472 13024 8488 13088
rect 8552 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8720 13088
rect 8400 12000 8720 13024
rect 8400 11936 8408 12000
rect 8472 11936 8488 12000
rect 8552 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8720 12000
rect 8400 10912 8720 11936
rect 8400 10848 8408 10912
rect 8472 10848 8488 10912
rect 8552 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8720 10912
rect 8400 9824 8720 10848
rect 8400 9760 8408 9824
rect 8472 9760 8488 9824
rect 8552 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8720 9824
rect 8400 9686 8720 9760
rect 8400 9450 8442 9686
rect 8678 9450 8720 9686
rect 8400 8736 8720 9450
rect 8400 8672 8408 8736
rect 8472 8672 8488 8736
rect 8552 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8720 8736
rect 8400 7648 8720 8672
rect 8400 7584 8408 7648
rect 8472 7584 8488 7648
rect 8552 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8720 7648
rect 8400 6560 8720 7584
rect 8400 6496 8408 6560
rect 8472 6496 8488 6560
rect 8552 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8720 6560
rect 8400 5472 8720 6496
rect 8400 5408 8408 5472
rect 8472 5408 8488 5472
rect 8552 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8720 5472
rect 8400 5198 8720 5408
rect 8400 4962 8442 5198
rect 8678 4962 8720 5198
rect 8400 4384 8720 4962
rect 8400 4320 8408 4384
rect 8472 4320 8488 4384
rect 8552 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8720 4384
rect 8400 3296 8720 4320
rect 8400 3232 8408 3296
rect 8472 3232 8488 3296
rect 8552 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8720 3296
rect 8400 2208 8720 3232
rect 8400 2144 8408 2208
rect 8472 2144 8488 2208
rect 8552 2144 8568 2208
rect 8632 2144 8648 2208
rect 8712 2144 8720 2208
rect 8400 2128 8720 2144
rect 12271 20160 12591 20176
rect 12271 20096 12279 20160
rect 12343 20096 12359 20160
rect 12423 20096 12439 20160
rect 12503 20096 12519 20160
rect 12583 20096 12591 20160
rect 12271 19072 12591 20096
rect 12271 19008 12279 19072
rect 12343 19008 12359 19072
rect 12423 19008 12439 19072
rect 12503 19008 12519 19072
rect 12583 19008 12591 19072
rect 12271 18002 12591 19008
rect 12271 17984 12313 18002
rect 12549 17984 12591 18002
rect 12271 17920 12279 17984
rect 12583 17920 12591 17984
rect 12271 17766 12313 17920
rect 12549 17766 12591 17920
rect 12271 16896 12591 17766
rect 12271 16832 12279 16896
rect 12343 16832 12359 16896
rect 12423 16832 12439 16896
rect 12503 16832 12519 16896
rect 12583 16832 12591 16896
rect 12271 15808 12591 16832
rect 12271 15744 12279 15808
rect 12343 15744 12359 15808
rect 12423 15744 12439 15808
rect 12503 15744 12519 15808
rect 12583 15744 12591 15808
rect 12271 14720 12591 15744
rect 12271 14656 12279 14720
rect 12343 14656 12359 14720
rect 12423 14656 12439 14720
rect 12503 14656 12519 14720
rect 12583 14656 12591 14720
rect 12271 13632 12591 14656
rect 12271 13568 12279 13632
rect 12343 13568 12359 13632
rect 12423 13568 12439 13632
rect 12503 13568 12519 13632
rect 12583 13568 12591 13632
rect 12271 13514 12591 13568
rect 12271 13278 12313 13514
rect 12549 13278 12591 13514
rect 12271 12544 12591 13278
rect 12271 12480 12279 12544
rect 12343 12480 12359 12544
rect 12423 12480 12439 12544
rect 12503 12480 12519 12544
rect 12583 12480 12591 12544
rect 12271 11456 12591 12480
rect 12271 11392 12279 11456
rect 12343 11392 12359 11456
rect 12423 11392 12439 11456
rect 12503 11392 12519 11456
rect 12583 11392 12591 11456
rect 12271 10368 12591 11392
rect 12271 10304 12279 10368
rect 12343 10304 12359 10368
rect 12423 10304 12439 10368
rect 12503 10304 12519 10368
rect 12583 10304 12591 10368
rect 12271 9280 12591 10304
rect 12271 9216 12279 9280
rect 12343 9216 12359 9280
rect 12423 9216 12439 9280
rect 12503 9216 12519 9280
rect 12583 9216 12591 9280
rect 12271 9026 12591 9216
rect 12271 8790 12313 9026
rect 12549 8790 12591 9026
rect 12271 8192 12591 8790
rect 12271 8128 12279 8192
rect 12343 8128 12359 8192
rect 12423 8128 12439 8192
rect 12503 8128 12519 8192
rect 12583 8128 12591 8192
rect 12271 7104 12591 8128
rect 12271 7040 12279 7104
rect 12343 7040 12359 7104
rect 12423 7040 12439 7104
rect 12503 7040 12519 7104
rect 12583 7040 12591 7104
rect 12271 6016 12591 7040
rect 12271 5952 12279 6016
rect 12343 5952 12359 6016
rect 12423 5952 12439 6016
rect 12503 5952 12519 6016
rect 12583 5952 12591 6016
rect 12271 4928 12591 5952
rect 12271 4864 12279 4928
rect 12343 4864 12359 4928
rect 12423 4864 12439 4928
rect 12503 4864 12519 4928
rect 12583 4864 12591 4928
rect 12271 4538 12591 4864
rect 12271 4302 12313 4538
rect 12549 4302 12591 4538
rect 12271 3840 12591 4302
rect 12271 3776 12279 3840
rect 12343 3776 12359 3840
rect 12423 3776 12439 3840
rect 12503 3776 12519 3840
rect 12583 3776 12591 3840
rect 12271 2752 12591 3776
rect 12271 2688 12279 2752
rect 12343 2688 12359 2752
rect 12423 2688 12439 2752
rect 12503 2688 12519 2752
rect 12583 2688 12591 2752
rect 12271 2128 12591 2688
rect 12931 19616 13251 20176
rect 12931 19552 12939 19616
rect 13003 19552 13019 19616
rect 13083 19552 13099 19616
rect 13163 19552 13179 19616
rect 13243 19552 13251 19616
rect 12931 18662 13251 19552
rect 12931 18528 12973 18662
rect 13209 18528 13251 18662
rect 12931 18464 12939 18528
rect 13243 18464 13251 18528
rect 12931 18426 12973 18464
rect 13209 18426 13251 18464
rect 12931 17440 13251 18426
rect 12931 17376 12939 17440
rect 13003 17376 13019 17440
rect 13083 17376 13099 17440
rect 13163 17376 13179 17440
rect 13243 17376 13251 17440
rect 12931 16352 13251 17376
rect 12931 16288 12939 16352
rect 13003 16288 13019 16352
rect 13083 16288 13099 16352
rect 13163 16288 13179 16352
rect 13243 16288 13251 16352
rect 12931 15264 13251 16288
rect 12931 15200 12939 15264
rect 13003 15200 13019 15264
rect 13083 15200 13099 15264
rect 13163 15200 13179 15264
rect 13243 15200 13251 15264
rect 12931 14176 13251 15200
rect 12931 14112 12939 14176
rect 13003 14174 13019 14176
rect 13083 14174 13099 14176
rect 13163 14174 13179 14176
rect 13243 14112 13251 14176
rect 12931 13938 12973 14112
rect 13209 13938 13251 14112
rect 12931 13088 13251 13938
rect 12931 13024 12939 13088
rect 13003 13024 13019 13088
rect 13083 13024 13099 13088
rect 13163 13024 13179 13088
rect 13243 13024 13251 13088
rect 12931 12000 13251 13024
rect 12931 11936 12939 12000
rect 13003 11936 13019 12000
rect 13083 11936 13099 12000
rect 13163 11936 13179 12000
rect 13243 11936 13251 12000
rect 12931 10912 13251 11936
rect 12931 10848 12939 10912
rect 13003 10848 13019 10912
rect 13083 10848 13099 10912
rect 13163 10848 13179 10912
rect 13243 10848 13251 10912
rect 12931 9824 13251 10848
rect 12931 9760 12939 9824
rect 13003 9760 13019 9824
rect 13083 9760 13099 9824
rect 13163 9760 13179 9824
rect 13243 9760 13251 9824
rect 12931 9686 13251 9760
rect 12931 9450 12973 9686
rect 13209 9450 13251 9686
rect 12931 8736 13251 9450
rect 12931 8672 12939 8736
rect 13003 8672 13019 8736
rect 13083 8672 13099 8736
rect 13163 8672 13179 8736
rect 13243 8672 13251 8736
rect 12931 7648 13251 8672
rect 12931 7584 12939 7648
rect 13003 7584 13019 7648
rect 13083 7584 13099 7648
rect 13163 7584 13179 7648
rect 13243 7584 13251 7648
rect 12931 6560 13251 7584
rect 12931 6496 12939 6560
rect 13003 6496 13019 6560
rect 13083 6496 13099 6560
rect 13163 6496 13179 6560
rect 13243 6496 13251 6560
rect 12931 5472 13251 6496
rect 12931 5408 12939 5472
rect 13003 5408 13019 5472
rect 13083 5408 13099 5472
rect 13163 5408 13179 5472
rect 13243 5408 13251 5472
rect 12931 5198 13251 5408
rect 12931 4962 12973 5198
rect 13209 4962 13251 5198
rect 12931 4384 13251 4962
rect 12931 4320 12939 4384
rect 13003 4320 13019 4384
rect 13083 4320 13099 4384
rect 13163 4320 13179 4384
rect 13243 4320 13251 4384
rect 12931 3296 13251 4320
rect 12931 3232 12939 3296
rect 13003 3232 13019 3296
rect 13083 3232 13099 3296
rect 13163 3232 13179 3296
rect 13243 3232 13251 3296
rect 12931 2208 13251 3232
rect 12931 2144 12939 2208
rect 13003 2144 13019 2208
rect 13083 2144 13099 2208
rect 13163 2144 13179 2208
rect 13243 2144 13251 2208
rect 12931 2128 13251 2144
rect 16802 20160 17122 20176
rect 16802 20096 16810 20160
rect 16874 20096 16890 20160
rect 16954 20096 16970 20160
rect 17034 20096 17050 20160
rect 17114 20096 17122 20160
rect 16802 19072 17122 20096
rect 16802 19008 16810 19072
rect 16874 19008 16890 19072
rect 16954 19008 16970 19072
rect 17034 19008 17050 19072
rect 17114 19008 17122 19072
rect 16802 18002 17122 19008
rect 16802 17984 16844 18002
rect 17080 17984 17122 18002
rect 16802 17920 16810 17984
rect 17114 17920 17122 17984
rect 16802 17766 16844 17920
rect 17080 17766 17122 17920
rect 16802 16896 17122 17766
rect 16802 16832 16810 16896
rect 16874 16832 16890 16896
rect 16954 16832 16970 16896
rect 17034 16832 17050 16896
rect 17114 16832 17122 16896
rect 16802 15808 17122 16832
rect 16802 15744 16810 15808
rect 16874 15744 16890 15808
rect 16954 15744 16970 15808
rect 17034 15744 17050 15808
rect 17114 15744 17122 15808
rect 16802 14720 17122 15744
rect 16802 14656 16810 14720
rect 16874 14656 16890 14720
rect 16954 14656 16970 14720
rect 17034 14656 17050 14720
rect 17114 14656 17122 14720
rect 16802 13632 17122 14656
rect 16802 13568 16810 13632
rect 16874 13568 16890 13632
rect 16954 13568 16970 13632
rect 17034 13568 17050 13632
rect 17114 13568 17122 13632
rect 16802 13514 17122 13568
rect 16802 13278 16844 13514
rect 17080 13278 17122 13514
rect 16802 12544 17122 13278
rect 16802 12480 16810 12544
rect 16874 12480 16890 12544
rect 16954 12480 16970 12544
rect 17034 12480 17050 12544
rect 17114 12480 17122 12544
rect 16802 11456 17122 12480
rect 16802 11392 16810 11456
rect 16874 11392 16890 11456
rect 16954 11392 16970 11456
rect 17034 11392 17050 11456
rect 17114 11392 17122 11456
rect 16802 10368 17122 11392
rect 16802 10304 16810 10368
rect 16874 10304 16890 10368
rect 16954 10304 16970 10368
rect 17034 10304 17050 10368
rect 17114 10304 17122 10368
rect 16802 9280 17122 10304
rect 16802 9216 16810 9280
rect 16874 9216 16890 9280
rect 16954 9216 16970 9280
rect 17034 9216 17050 9280
rect 17114 9216 17122 9280
rect 16802 9026 17122 9216
rect 16802 8790 16844 9026
rect 17080 8790 17122 9026
rect 16802 8192 17122 8790
rect 16802 8128 16810 8192
rect 16874 8128 16890 8192
rect 16954 8128 16970 8192
rect 17034 8128 17050 8192
rect 17114 8128 17122 8192
rect 16802 7104 17122 8128
rect 16802 7040 16810 7104
rect 16874 7040 16890 7104
rect 16954 7040 16970 7104
rect 17034 7040 17050 7104
rect 17114 7040 17122 7104
rect 16802 6016 17122 7040
rect 16802 5952 16810 6016
rect 16874 5952 16890 6016
rect 16954 5952 16970 6016
rect 17034 5952 17050 6016
rect 17114 5952 17122 6016
rect 16802 4928 17122 5952
rect 16802 4864 16810 4928
rect 16874 4864 16890 4928
rect 16954 4864 16970 4928
rect 17034 4864 17050 4928
rect 17114 4864 17122 4928
rect 16802 4538 17122 4864
rect 16802 4302 16844 4538
rect 17080 4302 17122 4538
rect 16802 3840 17122 4302
rect 16802 3776 16810 3840
rect 16874 3776 16890 3840
rect 16954 3776 16970 3840
rect 17034 3776 17050 3840
rect 17114 3776 17122 3840
rect 16802 2752 17122 3776
rect 16802 2688 16810 2752
rect 16874 2688 16890 2752
rect 16954 2688 16970 2752
rect 17034 2688 17050 2752
rect 17114 2688 17122 2752
rect 16802 2128 17122 2688
rect 17462 19616 17782 20176
rect 17462 19552 17470 19616
rect 17534 19552 17550 19616
rect 17614 19552 17630 19616
rect 17694 19552 17710 19616
rect 17774 19552 17782 19616
rect 17462 18662 17782 19552
rect 17462 18528 17504 18662
rect 17740 18528 17782 18662
rect 17462 18464 17470 18528
rect 17774 18464 17782 18528
rect 17462 18426 17504 18464
rect 17740 18426 17782 18464
rect 17462 17440 17782 18426
rect 17462 17376 17470 17440
rect 17534 17376 17550 17440
rect 17614 17376 17630 17440
rect 17694 17376 17710 17440
rect 17774 17376 17782 17440
rect 17462 16352 17782 17376
rect 17462 16288 17470 16352
rect 17534 16288 17550 16352
rect 17614 16288 17630 16352
rect 17694 16288 17710 16352
rect 17774 16288 17782 16352
rect 17462 15264 17782 16288
rect 17462 15200 17470 15264
rect 17534 15200 17550 15264
rect 17614 15200 17630 15264
rect 17694 15200 17710 15264
rect 17774 15200 17782 15264
rect 17462 14176 17782 15200
rect 17462 14112 17470 14176
rect 17534 14174 17550 14176
rect 17614 14174 17630 14176
rect 17694 14174 17710 14176
rect 17774 14112 17782 14176
rect 17462 13938 17504 14112
rect 17740 13938 17782 14112
rect 17462 13088 17782 13938
rect 17462 13024 17470 13088
rect 17534 13024 17550 13088
rect 17614 13024 17630 13088
rect 17694 13024 17710 13088
rect 17774 13024 17782 13088
rect 17462 12000 17782 13024
rect 17462 11936 17470 12000
rect 17534 11936 17550 12000
rect 17614 11936 17630 12000
rect 17694 11936 17710 12000
rect 17774 11936 17782 12000
rect 17462 10912 17782 11936
rect 17462 10848 17470 10912
rect 17534 10848 17550 10912
rect 17614 10848 17630 10912
rect 17694 10848 17710 10912
rect 17774 10848 17782 10912
rect 17462 9824 17782 10848
rect 17462 9760 17470 9824
rect 17534 9760 17550 9824
rect 17614 9760 17630 9824
rect 17694 9760 17710 9824
rect 17774 9760 17782 9824
rect 17462 9686 17782 9760
rect 17462 9450 17504 9686
rect 17740 9450 17782 9686
rect 17462 8736 17782 9450
rect 17462 8672 17470 8736
rect 17534 8672 17550 8736
rect 17614 8672 17630 8736
rect 17694 8672 17710 8736
rect 17774 8672 17782 8736
rect 17462 7648 17782 8672
rect 17462 7584 17470 7648
rect 17534 7584 17550 7648
rect 17614 7584 17630 7648
rect 17694 7584 17710 7648
rect 17774 7584 17782 7648
rect 17462 6560 17782 7584
rect 17462 6496 17470 6560
rect 17534 6496 17550 6560
rect 17614 6496 17630 6560
rect 17694 6496 17710 6560
rect 17774 6496 17782 6560
rect 17462 5472 17782 6496
rect 17462 5408 17470 5472
rect 17534 5408 17550 5472
rect 17614 5408 17630 5472
rect 17694 5408 17710 5472
rect 17774 5408 17782 5472
rect 17462 5198 17782 5408
rect 17462 4962 17504 5198
rect 17740 4962 17782 5198
rect 17462 4384 17782 4962
rect 17462 4320 17470 4384
rect 17534 4320 17550 4384
rect 17614 4320 17630 4384
rect 17694 4320 17710 4384
rect 17774 4320 17782 4384
rect 17462 3296 17782 4320
rect 17462 3232 17470 3296
rect 17534 3232 17550 3296
rect 17614 3232 17630 3296
rect 17694 3232 17710 3296
rect 17774 3232 17782 3296
rect 17462 2208 17782 3232
rect 17462 2144 17470 2208
rect 17534 2144 17550 2208
rect 17614 2144 17630 2208
rect 17694 2144 17710 2208
rect 17774 2144 17782 2208
rect 17462 2128 17782 2144
<< via4 >>
rect 3251 17984 3487 18002
rect 3251 17920 3281 17984
rect 3281 17920 3297 17984
rect 3297 17920 3361 17984
rect 3361 17920 3377 17984
rect 3377 17920 3441 17984
rect 3441 17920 3457 17984
rect 3457 17920 3487 17984
rect 3251 17766 3487 17920
rect 3251 13278 3487 13514
rect 3251 8790 3487 9026
rect 3251 4302 3487 4538
rect 3911 18528 4147 18662
rect 3911 18464 3941 18528
rect 3941 18464 3957 18528
rect 3957 18464 4021 18528
rect 4021 18464 4037 18528
rect 4037 18464 4101 18528
rect 4101 18464 4117 18528
rect 4117 18464 4147 18528
rect 3911 18426 4147 18464
rect 3911 14112 3941 14174
rect 3941 14112 3957 14174
rect 3957 14112 4021 14174
rect 4021 14112 4037 14174
rect 4037 14112 4101 14174
rect 4101 14112 4117 14174
rect 4117 14112 4147 14174
rect 3911 13938 4147 14112
rect 7782 17984 8018 18002
rect 7782 17920 7812 17984
rect 7812 17920 7828 17984
rect 7828 17920 7892 17984
rect 7892 17920 7908 17984
rect 7908 17920 7972 17984
rect 7972 17920 7988 17984
rect 7988 17920 8018 17984
rect 7782 17766 8018 17920
rect 7782 13278 8018 13514
rect 3911 9450 4147 9686
rect 7782 8790 8018 9026
rect 3911 4962 4147 5198
rect 7782 4302 8018 4538
rect 8442 18528 8678 18662
rect 8442 18464 8472 18528
rect 8472 18464 8488 18528
rect 8488 18464 8552 18528
rect 8552 18464 8568 18528
rect 8568 18464 8632 18528
rect 8632 18464 8648 18528
rect 8648 18464 8678 18528
rect 8442 18426 8678 18464
rect 8442 14112 8472 14174
rect 8472 14112 8488 14174
rect 8488 14112 8552 14174
rect 8552 14112 8568 14174
rect 8568 14112 8632 14174
rect 8632 14112 8648 14174
rect 8648 14112 8678 14174
rect 8442 13938 8678 14112
rect 8442 9450 8678 9686
rect 8442 4962 8678 5198
rect 12313 17984 12549 18002
rect 12313 17920 12343 17984
rect 12343 17920 12359 17984
rect 12359 17920 12423 17984
rect 12423 17920 12439 17984
rect 12439 17920 12503 17984
rect 12503 17920 12519 17984
rect 12519 17920 12549 17984
rect 12313 17766 12549 17920
rect 12313 13278 12549 13514
rect 12313 8790 12549 9026
rect 12313 4302 12549 4538
rect 12973 18528 13209 18662
rect 12973 18464 13003 18528
rect 13003 18464 13019 18528
rect 13019 18464 13083 18528
rect 13083 18464 13099 18528
rect 13099 18464 13163 18528
rect 13163 18464 13179 18528
rect 13179 18464 13209 18528
rect 12973 18426 13209 18464
rect 12973 14112 13003 14174
rect 13003 14112 13019 14174
rect 13019 14112 13083 14174
rect 13083 14112 13099 14174
rect 13099 14112 13163 14174
rect 13163 14112 13179 14174
rect 13179 14112 13209 14174
rect 12973 13938 13209 14112
rect 12973 9450 13209 9686
rect 12973 4962 13209 5198
rect 16844 17984 17080 18002
rect 16844 17920 16874 17984
rect 16874 17920 16890 17984
rect 16890 17920 16954 17984
rect 16954 17920 16970 17984
rect 16970 17920 17034 17984
rect 17034 17920 17050 17984
rect 17050 17920 17080 17984
rect 16844 17766 17080 17920
rect 16844 13278 17080 13514
rect 16844 8790 17080 9026
rect 16844 4302 17080 4538
rect 17504 18528 17740 18662
rect 17504 18464 17534 18528
rect 17534 18464 17550 18528
rect 17550 18464 17614 18528
rect 17614 18464 17630 18528
rect 17630 18464 17694 18528
rect 17694 18464 17710 18528
rect 17710 18464 17740 18528
rect 17504 18426 17740 18464
rect 17504 14112 17534 14174
rect 17534 14112 17550 14174
rect 17550 14112 17614 14174
rect 17614 14112 17630 14174
rect 17630 14112 17694 14174
rect 17694 14112 17710 14174
rect 17710 14112 17740 14174
rect 17504 13938 17740 14112
rect 17504 9450 17740 9686
rect 17504 4962 17740 5198
<< metal5 >>
rect 1056 18662 19276 18704
rect 1056 18426 3911 18662
rect 4147 18426 8442 18662
rect 8678 18426 12973 18662
rect 13209 18426 17504 18662
rect 17740 18426 19276 18662
rect 1056 18384 19276 18426
rect 1056 18002 19276 18044
rect 1056 17766 3251 18002
rect 3487 17766 7782 18002
rect 8018 17766 12313 18002
rect 12549 17766 16844 18002
rect 17080 17766 19276 18002
rect 1056 17724 19276 17766
rect 1056 14174 19276 14216
rect 1056 13938 3911 14174
rect 4147 13938 8442 14174
rect 8678 13938 12973 14174
rect 13209 13938 17504 14174
rect 17740 13938 19276 14174
rect 1056 13896 19276 13938
rect 1056 13514 19276 13556
rect 1056 13278 3251 13514
rect 3487 13278 7782 13514
rect 8018 13278 12313 13514
rect 12549 13278 16844 13514
rect 17080 13278 19276 13514
rect 1056 13236 19276 13278
rect 1056 9686 19276 9728
rect 1056 9450 3911 9686
rect 4147 9450 8442 9686
rect 8678 9450 12973 9686
rect 13209 9450 17504 9686
rect 17740 9450 19276 9686
rect 1056 9408 19276 9450
rect 1056 9026 19276 9068
rect 1056 8790 3251 9026
rect 3487 8790 7782 9026
rect 8018 8790 12313 9026
rect 12549 8790 16844 9026
rect 17080 8790 19276 9026
rect 1056 8748 19276 8790
rect 1056 5198 19276 5240
rect 1056 4962 3911 5198
rect 4147 4962 8442 5198
rect 8678 4962 12973 5198
rect 13209 4962 17504 5198
rect 17740 4962 19276 5198
rect 1056 4920 19276 4962
rect 1056 4538 19276 4580
rect 1056 4302 3251 4538
rect 3487 4302 7782 4538
rect 8018 4302 12313 4538
rect 12549 4302 16844 4538
rect 17080 4302 19276 4538
rect 1056 4260 19276 4302
use sky130_fd_sc_hd__clkbuf_4  _206_
timestamp 0
transform 1 0 1748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _207_
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _208_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _209_
timestamp 0
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _210_
timestamp 0
transform -1 0 3588 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _211_
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp 0
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _213_
timestamp 0
transform -1 0 3864 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _214_
timestamp 0
transform 1 0 9752 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _215_
timestamp 0
transform 1 0 10304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 0
transform 1 0 9292 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _218_
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _219_
timestamp 0
transform -1 0 9384 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _220_
timestamp 0
transform -1 0 5612 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _221_
timestamp 0
transform -1 0 4784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _222_
timestamp 0
transform 1 0 4324 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _223_
timestamp 0
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 0
transform -1 0 7452 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _225_
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _226_
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _227_
timestamp 0
transform -1 0 8464 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _228_
timestamp 0
transform 1 0 1840 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _229_
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _230_
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 0
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _232_
timestamp 0
transform 1 0 3312 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _233_
timestamp 0
transform -1 0 4140 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _234_
timestamp 0
transform -1 0 3036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _235_
timestamp 0
transform 1 0 2116 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _236_
timestamp 0
transform -1 0 3496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _237_
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _238_
timestamp 0
transform -1 0 5244 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _239_
timestamp 0
transform -1 0 6072 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _240_
timestamp 0
transform 1 0 4232 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 0
transform -1 0 4140 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _242_
timestamp 0
transform 1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _243_
timestamp 0
transform -1 0 2852 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 0
transform -1 0 3680 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _245_
timestamp 0
transform 1 0 2300 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _246_
timestamp 0
transform 1 0 4508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _247_
timestamp 0
transform 1 0 2944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _248_
timestamp 0
transform 1 0 2208 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _249_
timestamp 0
transform -1 0 3864 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _250_
timestamp 0
transform -1 0 5060 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _251_
timestamp 0
transform 1 0 2760 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp 0
transform -1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _253_
timestamp 0
transform -1 0 3128 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _254_
timestamp 0
transform -1 0 6992 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _255_
timestamp 0
transform -1 0 7820 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _256_
timestamp 0
transform 1 0 5152 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _257_
timestamp 0
transform -1 0 4968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _258_
timestamp 0
transform -1 0 4416 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _259_
timestamp 0
transform -1 0 5336 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _260_
timestamp 0
transform -1 0 5796 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _261_
timestamp 0
transform 1 0 4600 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 0
transform -1 0 6164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _263_
timestamp 0
transform 1 0 5244 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _264_
timestamp 0
transform 1 0 12144 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _265_
timestamp 0
transform -1 0 7728 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _266_
timestamp 0
transform -1 0 7912 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _267_
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _268_
timestamp 0
transform -1 0 7268 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _269_
timestamp 0
transform -1 0 6992 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _270_
timestamp 0
transform -1 0 7176 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _271_
timestamp 0
transform -1 0 8004 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _272_
timestamp 0
transform 1 0 6440 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _273_
timestamp 0
transform -1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _274_
timestamp 0
transform -1 0 6992 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _275_
timestamp 0
transform -1 0 10396 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 0
transform -1 0 9660 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _277_
timestamp 0
transform 1 0 8924 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _278_
timestamp 0
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _279_
timestamp 0
transform 1 0 8188 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _280_
timestamp 0
transform -1 0 8648 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _281_
timestamp 0
transform -1 0 8740 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _282_
timestamp 0
transform 1 0 7360 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _283_
timestamp 0
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _284_
timestamp 0
transform 1 0 7912 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _285_
timestamp 0
transform -1 0 9476 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _286_
timestamp 0
transform -1 0 10120 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _287_
timestamp 0
transform 1 0 8096 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 0
transform -1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _289_
timestamp 0
transform 1 0 8280 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _290_
timestamp 0
transform -1 0 12604 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 0
transform -1 0 13064 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _292_
timestamp 0
transform 1 0 10028 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 0
transform -1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _294_
timestamp 0
transform 1 0 9752 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _295_
timestamp 0
transform -1 0 13156 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp 0
transform -1 0 11960 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _297_
timestamp 0
transform 1 0 10488 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _298_
timestamp 0
transform -1 0 15824 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _299_
timestamp 0
transform 1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _300_
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _301_
timestamp 0
transform -1 0 11132 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _302_
timestamp 0
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _303_
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _304_
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _305_
timestamp 0
transform 1 0 10488 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _306_
timestamp 0
transform -1 0 13984 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _307_
timestamp 0
transform -1 0 14536 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 0
transform 1 0 12236 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _309_
timestamp 0
transform -1 0 11408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _310_
timestamp 0
transform -1 0 11316 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _311_
timestamp 0
transform -1 0 14444 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _312_
timestamp 0
transform -1 0 13248 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _313_
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _314_
timestamp 0
transform 1 0 12880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _315_
timestamp 0
transform 1 0 12328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _316_
timestamp 0
transform 1 0 11500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _317_
timestamp 0
transform -1 0 14720 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _318_
timestamp 0
transform -1 0 15732 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _319_
timestamp 0
transform 1 0 13064 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _320_
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _321_
timestamp 0
transform -1 0 13800 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _322_
timestamp 0
transform -1 0 14720 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp 0
transform -1 0 14628 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _324_
timestamp 0
transform 1 0 13064 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _325_
timestamp 0
transform -1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _326_
timestamp 0
transform 1 0 13156 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _327_
timestamp 0
transform -1 0 18216 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 0
transform -1 0 18952 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _329_
timestamp 0
transform 1 0 16652 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 0
transform -1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _331_
timestamp 0
transform -1 0 15640 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _332_
timestamp 0
transform -1 0 18768 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _333_
timestamp 0
transform -1 0 18124 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _334_
timestamp 0
transform -1 0 16284 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 0
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _336_
timestamp 0
transform 1 0 15732 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _337_
timestamp 0
transform -1 0 17756 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _338_
timestamp 0
transform -1 0 18400 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _339_
timestamp 0
transform 1 0 15640 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _340_
timestamp 0
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _341_
timestamp 0
transform 1 0 16652 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _342_
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 0
transform -1 0 16192 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _344_
timestamp 0
transform 1 0 15272 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _345_
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _346_
timestamp 0
transform -1 0 18308 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _347_
timestamp 0
transform -1 0 18492 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _348_
timestamp 0
transform -1 0 18952 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _349_
timestamp 0
transform 1 0 16560 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _350_
timestamp 0
transform -1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _351_
timestamp 0
transform -1 0 15456 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _352_
timestamp 0
transform -1 0 18216 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _353_
timestamp 0
transform -1 0 18952 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _354_
timestamp 0
transform -1 0 16560 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 0
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _356_
timestamp 0
transform 1 0 15640 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _357_
timestamp 0
transform -1 0 16468 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _358_
timestamp 0
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _359_
timestamp 0
transform 1 0 15824 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _360_
timestamp 0
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _361_
timestamp 0
transform 1 0 16560 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _362_
timestamp 0
transform 1 0 14720 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 0
transform 1 0 13524 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _364_
timestamp 0
transform 1 0 14812 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _365_
timestamp 0
transform -1 0 15732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _366_
timestamp 0
transform -1 0 15548 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 0
transform -1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _368_
timestamp 0
transform -1 0 13432 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _369_
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 0
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _371_
timestamp 0
transform 1 0 12328 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _372_
timestamp 0
transform -1 0 15456 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _373_
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 0
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 0
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 0
transform 1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 0
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 0
transform -1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 0
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 0
transform 1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 0
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 0
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _384_
timestamp 0
transform -1 0 6900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 0
transform 1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 0
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 0
transform 1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 0
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 0
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 0
transform -1 0 3680 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 0
transform -1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 0
transform -1 0 6072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 0
transform -1 0 1840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _395_
timestamp 0
transform -1 0 6256 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 0
transform -1 0 4692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 0
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 0
transform -1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 0
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 0
transform 1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 0
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 0
transform 1 0 9016 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _406_
timestamp 0
transform 1 0 9016 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 0
transform -1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 0
transform -1 0 10028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 0
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 0
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 0
transform 1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 0
transform 1 0 11868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 0
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 0
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 0
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _417_
timestamp 0
transform 1 0 14720 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 0
transform -1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 0
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 0
transform -1 0 13984 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 0
transform -1 0 14996 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 0
transform -1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 0
transform -1 0 15732 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 0
transform 1 0 17296 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 0
transform -1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 0
transform 1 0 17296 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 0
transform 1 0 17572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _428_
timestamp 0
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 0
transform 1 0 15824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 0
transform 1 0 18400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 0
transform -1 0 15548 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 0
transform -1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 0
transform 1 0 17572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 0
transform -1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 0
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 0
transform 1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 0
transform 1 0 15548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 0
transform -1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 0
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 0
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 0
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 0
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _443_
timestamp 0
transform 1 0 1748 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _444_
timestamp 0
transform -1 0 3220 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 0
transform 1 0 7912 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp 0
transform 1 0 8924 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _447_
timestamp 0
transform 1 0 5612 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _448_
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _449_
timestamp 0
transform 1 0 4140 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _450_
timestamp 0
transform 1 0 7084 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _451_
timestamp 0
transform -1 0 3220 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _452_
timestamp 0
transform 1 0 4232 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _453_
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _454_
timestamp 0
transform -1 0 3220 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _455_
timestamp 0
transform 1 0 3864 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _456_
timestamp 0
transform 1 0 4140 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _457_
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _458_
timestamp 0
transform 1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 0
transform 1 0 1840 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 0
transform -1 0 3220 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _461_
timestamp 0
transform 1 0 4416 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _462_
timestamp 0
transform -1 0 3220 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp 0
transform 1 0 5428 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 0
transform 1 0 7912 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 0
transform -1 0 9752 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 0
transform 1 0 6440 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 0
transform 1 0 8280 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _473_
timestamp 0
transform 1 0 6992 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _474_
timestamp 0
transform -1 0 10764 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 0
transform 1 0 10120 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 0
transform 1 0 10304 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _479_
timestamp 0
transform 1 0 9292 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _480_
timestamp 0
transform 1 0 10764 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _481_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 0
transform 1 0 9108 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 0
transform 1 0 11960 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 0
transform -1 0 14720 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _485_
timestamp 0
transform 1 0 12144 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _486_
timestamp 0
transform 1 0 12880 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _487_
timestamp 0
transform 1 0 12328 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 0
transform 1 0 13616 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 0
transform 1 0 14904 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 0
transform 1 0 16744 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 0
transform 1 0 14996 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 0
transform 1 0 17112 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 0
transform 1 0 14260 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 0
transform 1 0 17112 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _498_
timestamp 0
transform 1 0 14352 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 0
transform 1 0 14536 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 0
transform 1 0 17112 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp 0
transform 1 0 11868 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 0
transform 1 0 14168 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _505_
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 0
transform 1 0 12236 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 11132 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 0
transform -1 0 3680 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 0
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 0
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 0
transform 1 0 5244 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 0
transform -1 0 12236 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 0
transform 1 0 13340 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 0
transform -1 0 12236 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 0
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_157
timestamp 0
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_193
timestamp 0
transform 1 0 18860 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_20
timestamp 0
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_32
timestamp 0
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_44
timestamp 0
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_156
timestamp 0
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_36
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_48
timestamp 0
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_52
timestamp 0
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_64
timestamp 0
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_76
timestamp 0
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_89
timestamp 0
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_93
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_105
timestamp 0
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_117
timestamp 0
transform 1 0 11868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_129
timestamp 0
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_135
timestamp 0
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_149
timestamp 0
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_154
timestamp 0
transform 1 0 15272 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_166
timestamp 0
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_178
timestamp 0
transform 1 0 17480 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_190
timestamp 0
transform 1 0 18584 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_21
timestamp 0
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_35
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_63
timestamp 0
transform 1 0 6900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_75
timestamp 0
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_120
timestamp 0
transform 1 0 12144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 0
transform 1 0 14076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_162
timestamp 0
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_9
timestamp 0
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 0
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_113
timestamp 0
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_134
timestamp 0
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_159
timestamp 0
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_167
timestamp 0
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_175
timestamp 0
transform 1 0 17204 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_183
timestamp 0
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_193
timestamp 0
transform 1 0 18860 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_30
timestamp 0
transform 1 0 3864 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_36
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_40
timestamp 0
transform 1 0 4784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_52
timestamp 0
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_96
timestamp 0
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_102
timestamp 0
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 0
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_128
timestamp 0
transform 1 0 12880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_140
timestamp 0
transform 1 0 13984 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 0
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_11
timestamp 0
transform 1 0 2116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_19
timestamp 0
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_35
timestamp 0
transform 1 0 4324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_45
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 0
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 0
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_88
timestamp 0
transform 1 0 9200 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_94
timestamp 0
transform 1 0 9752 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_106
timestamp 0
transform 1 0 10856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_112
timestamp 0
transform 1 0 11408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_122
timestamp 0
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_126
timestamp 0
transform 1 0 12696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_130
timestamp 0
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 0
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_167
timestamp 0
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_184
timestamp 0
transform 1 0 18032 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_192
timestamp 0
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_23
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_31
timestamp 0
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 0
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 0
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_155
timestamp 0
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_172
timestamp 0
transform 1 0 16928 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_184
timestamp 0
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_188
timestamp 0
transform 1 0 18400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_89
timestamp 0
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_124
timestamp 0
transform 1 0 12512 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_132
timestamp 0
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_162
timestamp 0
transform 1 0 16008 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_174
timestamp 0
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_22
timestamp 0
transform 1 0 3128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_66
timestamp 0
transform 1 0 7176 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_78
timestamp 0
transform 1 0 8280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_86
timestamp 0
transform 1 0 9016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_107
timestamp 0
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_159
timestamp 0
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_189
timestamp 0
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_193
timestamp 0
transform 1 0 18860 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 0
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 0
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_92
timestamp 0
transform 1 0 9568 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_111
timestamp 0
transform 1 0 11316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_123
timestamp 0
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_149
timestamp 0
transform 1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp 0
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_189
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_193
timestamp 0
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_9
timestamp 0
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_20
timestamp 0
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_32
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_40
timestamp 0
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_45
timestamp 0
transform 1 0 5244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_49
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_94
timestamp 0
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_106
timestamp 0
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_154
timestamp 0
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 0
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_192
timestamp 0
transform 1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 0
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_57
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 0
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_88
timestamp 0
transform 1 0 9200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_100
timestamp 0
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_119
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_126
timestamp 0
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_130
timestamp 0
transform 1 0 13064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_167
timestamp 0
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_175
timestamp 0
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_189
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_193
timestamp 0
transform 1 0 18860 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_47
timestamp 0
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_63
timestamp 0
transform 1 0 6900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_75
timestamp 0
transform 1 0 8004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_87
timestamp 0
transform 1 0 9108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_118
timestamp 0
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_129
timestamp 0
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_141
timestamp 0
transform 1 0 14076 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_159
timestamp 0
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_21
timestamp 0
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_67
timestamp 0
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 0
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_108
timestamp 0
transform 1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_112
timestamp 0
transform 1 0 11408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_131
timestamp 0
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 0
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_185
timestamp 0
transform 1 0 18124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_7
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_33
timestamp 0
transform 1 0 4140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_84
timestamp 0
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_95
timestamp 0
transform 1 0 9844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 0
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_117
timestamp 0
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_145
timestamp 0
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_153
timestamp 0
transform 1 0 15180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_157
timestamp 0
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 0
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_176
timestamp 0
transform 1 0 17296 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_188
timestamp 0
transform 1 0 18400 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_23
timestamp 0
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_61
timestamp 0
transform 1 0 6716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_112
timestamp 0
transform 1 0 11408 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_124
timestamp 0
transform 1 0 12512 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_163
timestamp 0
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_190
timestamp 0
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_101
timestamp 0
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 0
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_118
timestamp 0
transform 1 0 11960 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_126
timestamp 0
transform 1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_153
timestamp 0
transform 1 0 15180 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp 0
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 0
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_32
timestamp 0
transform 1 0 4048 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_72
timestamp 0
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_101
timestamp 0
transform 1 0 10396 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_125
timestamp 0
transform 1 0 12604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 0
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_176
timestamp 0
transform 1 0 17296 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_188
timestamp 0
transform 1 0 18400 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_11
timestamp 0
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_19
timestamp 0
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_31
timestamp 0
transform 1 0 3956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_43
timestamp 0
transform 1 0 5060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_77
timestamp 0
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_98
timestamp 0
transform 1 0 10120 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 0
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_118
timestamp 0
transform 1 0 11960 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_126
timestamp 0
transform 1 0 12696 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_151
timestamp 0
transform 1 0 14996 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_157
timestamp 0
transform 1 0 15548 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 0
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_191
timestamp 0
transform 1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_9
timestamp 0
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_23
timestamp 0
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_52
timestamp 0
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_56
timestamp 0
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 0
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_89
timestamp 0
transform 1 0 9292 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_115
timestamp 0
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 0
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_149
timestamp 0
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_171
timestamp 0
transform 1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_28
timestamp 0
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_40
timestamp 0
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 0
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_67
timestamp 0
transform 1 0 7268 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_79
timestamp 0
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_91
timestamp 0
transform 1 0 9476 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_99
timestamp 0
transform 1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 0
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_121
timestamp 0
transform 1 0 12236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 0
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_140
timestamp 0
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_148
timestamp 0
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 0
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_173
timestamp 0
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_11
timestamp 0
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_19
timestamp 0
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_37
timestamp 0
transform 1 0 4508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_49
timestamp 0
transform 1 0 5612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_61
timestamp 0
transform 1 0 6716 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_70
timestamp 0
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_93
timestamp 0
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_105
timestamp 0
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_111
timestamp 0
transform 1 0 11316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_145
timestamp 0
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_159
timestamp 0
transform 1 0 15732 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_171
timestamp 0
transform 1 0 16836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_183
timestamp 0
transform 1 0 17940 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_191
timestamp 0
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_13
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_25
timestamp 0
transform 1 0 3404 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_33
timestamp 0
transform 1 0 4140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_83
timestamp 0
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_133
timestamp 0
transform 1 0 13340 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_140
timestamp 0
transform 1 0 13984 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_152
timestamp 0
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 0
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_175
timestamp 0
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_179
timestamp 0
transform 1 0 17572 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_192
timestamp 0
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 0
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_57
timestamp 0
transform 1 0 6348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_61
timestamp 0
transform 1 0 6716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_67
timestamp 0
transform 1 0 7268 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_75
timestamp 0
transform 1 0 8004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_93
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_157
timestamp 0
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_185
timestamp 0
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_6
timestamp 0
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_10
timestamp 0
transform 1 0 2024 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_14
timestamp 0
transform 1 0 2392 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_25
timestamp 0
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_37
timestamp 0
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_82
timestamp 0
transform 1 0 8648 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_94
timestamp 0
transform 1 0 9752 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_106
timestamp 0
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_117
timestamp 0
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_130
timestamp 0
transform 1 0 13064 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 0
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_177
timestamp 0
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_182
timestamp 0
transform 1 0 17848 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_67
timestamp 0
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 0
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_118
timestamp 0
transform 1 0 11960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_122
timestamp 0
transform 1 0 12328 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 0
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_157
timestamp 0
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_161
timestamp 0
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_169
timestamp 0
transform 1 0 16652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_190
timestamp 0
transform 1 0 18584 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_30
timestamp 0
transform 1 0 3864 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_38
timestamp 0
transform 1 0 4600 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_42
timestamp 0
transform 1 0 4968 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_50
timestamp 0
transform 1 0 5704 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 0
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_64
timestamp 0
transform 1 0 6992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_76
timestamp 0
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_88
timestamp 0
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_131
timestamp 0
transform 1 0 13156 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_135
timestamp 0
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_147
timestamp 0
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_158
timestamp 0
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 0
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_43
timestamp 0
transform 1 0 5060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_51
timestamp 0
transform 1 0 5796 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_73
timestamp 0
transform 1 0 7820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_98
timestamp 0
transform 1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_120
timestamp 0
transform 1 0 12144 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_128
timestamp 0
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 0
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_148
timestamp 0
transform 1 0 14720 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_173
timestamp 0
transform 1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_28
timestamp 0
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 0
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_91
timestamp 0
transform 1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_104
timestamp 0
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_116
timestamp 0
transform 1 0 11776 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_142
timestamp 0
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_152
timestamp 0
transform 1 0 15088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_156
timestamp 0
transform 1 0 15456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 0
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_189
timestamp 0
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_193
timestamp 0
transform 1 0 18860 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_9
timestamp 0
transform 1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_21
timestamp 0
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_33
timestamp 0
transform 1 0 4140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_39
timestamp 0
transform 1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_45
timestamp 0
transform 1 0 5244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_51
timestamp 0
transform 1 0 5796 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_55
timestamp 0
transform 1 0 6164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_63
timestamp 0
transform 1 0 6900 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_69
timestamp 0
transform 1 0 7452 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_75
timestamp 0
transform 1 0 8004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 0
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_88
timestamp 0
transform 1 0 9200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_93
timestamp 0
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_99
timestamp 0
transform 1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_105
timestamp 0
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_111
timestamp 0
transform 1 0 11316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_113
timestamp 0
transform 1 0 11500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_117
timestamp 0
transform 1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_123
timestamp 0
transform 1 0 12420 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_129
timestamp 0
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_159
timestamp 0
transform 1 0 15732 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_185
timestamp 0
transform 1 0 18124 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_189
timestamp 0
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 8556 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 8924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 8188 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 8832 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform 1 0 11592 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 12880 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 5152 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 3496 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform 1 0 14352 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 11408 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 8556 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 7728 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 16284 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform -1 0 8832 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform 1 0 16928 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform -1 0 12512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 12236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 7912 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 13984 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 13340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 0
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 0
transform -1 0 5612 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 0
transform -1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 0
transform -1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 0
transform 1 0 13984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 0
transform 1 0 3864 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 0
transform -1 0 18032 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 0
transform -1 0 17296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 0
transform 1 0 12420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 0
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 0
transform 1 0 6624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 0
transform -1 0 6624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 0
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 0
transform -1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 0
transform -1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 0
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 0
transform 1 0 17204 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 0
transform 1 0 14536 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 0
transform -1 0 18952 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 0
transform -1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 0
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 0
transform 1 0 18216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 0
transform 1 0 11316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 0
transform -1 0 14904 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform -1 0 7452 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform -1 0 8004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 8280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform -1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 9384 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform 1 0 10488 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform 1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform 1 0 11592 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 0
transform 1 0 12144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 0
transform 1 0 2208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 0
transform 1 0 12696 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform 1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform 1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 0
transform 1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 0
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 0
transform -1 0 17572 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 0
transform -1 0 17848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 0
transform -1 0 18124 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 0
transform 1 0 2760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 0
transform -1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 0
transform -1 0 18952 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 0
transform 1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 0
transform -1 0 4140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 0
transform 1 0 4416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 0
transform -1 0 5244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 0
transform -1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 0
transform -1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 0
transform -1 0 6900 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 0
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 19228 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 19228 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 19228 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 19228 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 19228 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 19228 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 19228 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 19228 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 6256 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 11408 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 16560 0 1 19584
box -38 -48 130 592
<< labels >>
rlabel metal1 s 10166 19584 10166 19584 4 VGND
rlabel metal1 s 10166 20128 10166 20128 4 VPWR
rlabel metal1 s 2300 4658 2300 4658 4 _000_
rlabel metal1 s 6624 13974 6624 13974 4 _001_
rlabel metal1 s 6532 8874 6532 8874 4 _002_
rlabel metal1 s 8602 12750 8602 12750 4 _003_
rlabel metal1 s 7084 16014 7084 16014 4 _004_
rlabel metal1 s 7728 18938 7728 18938 4 _005_
rlabel metal1 s 10258 17714 10258 17714 4 _006_
rlabel metal1 s 10343 14586 10343 14586 4 _007_
rlabel metal1 s 9614 10744 9614 10744 4 _008_
rlabel metal1 s 11822 8568 11822 8568 4 _009_
rlabel metal1 s 12236 11254 12236 11254 4 _010_
rlabel metal1 s 5750 5746 5750 5746 4 _011_
rlabel metal1 s 12788 15130 12788 15130 4 _012_
rlabel metal1 s 12880 18938 12880 18938 4 _013_
rlabel metal1 s 16974 19448 16974 19448 4 _014_
rlabel metal1 s 16606 16456 16606 16456 4 _015_
rlabel metal1 s 15502 14042 15502 14042 4 _016_
rlabel metal1 s 14950 12274 14950 12274 4 _017_
rlabel metal2 s 16606 10370 16606 10370 4 _018_
rlabel metal1 s 16744 8398 16744 8398 4 _019_
rlabel metal1 s 15364 6222 15364 6222 4 _020_
rlabel metal1 s 13662 7344 13662 7344 4 _021_
rlabel metal1 s 4462 7480 4462 7480 4 _022_
rlabel metal1 s 10757 5882 10757 5882 4 _023_
rlabel metal1 s 2714 8296 2714 8296 4 _024_
rlabel metal1 s 2162 11832 2162 11832 4 _025_
rlabel metal2 s 4278 12002 4278 12002 4 _026_
rlabel metal1 s 2024 14586 2024 14586 4 _027_
rlabel metal1 s 2162 18632 2162 18632 4 _028_
rlabel metal1 s 4968 18938 4968 18938 4 _029_
rlabel metal1 s 4370 16626 4370 16626 4 _030_
rlabel metal1 s 9246 5304 9246 5304 4 _031_
rlabel metal1 s 9016 7310 9016 7310 4 _032_
rlabel metal2 s 2806 4386 2806 4386 4 _033_
rlabel metal1 s 2300 5882 2300 5882 4 _034_
rlabel metal1 s 9016 6970 9016 6970 4 _035_
rlabel metal1 s 9614 4794 9614 4794 4 _036_
rlabel metal1 s 6854 5338 6854 5338 4 _037_
rlabel metal2 s 5750 5032 5750 5032 4 _038_
rlabel metal1 s 5336 6766 5336 6766 4 _039_
rlabel metal2 s 9522 6120 9522 6120 4 _040_
rlabel metal1 s 2300 6970 2300 6970 4 _041_
rlabel metal1 s 5014 8058 5014 8058 4 _042_
rlabel metal2 s 1978 12002 1978 12002 4 _043_
rlabel metal2 s 2162 9826 2162 9826 4 _044_
rlabel metal1 s 5987 12138 5987 12138 4 _045_
rlabel metal1 s 5244 10438 5244 10438 4 _046_
rlabel metal2 s 2162 14790 2162 14790 4 _047_
rlabel metal1 s 5053 12886 5053 12886 4 _048_
rlabel metal2 s 2622 18938 2622 18938 4 _049_
rlabel metal2 s 2254 16728 2254 16728 4 _050_
rlabel metal1 s 5888 18394 5888 18394 4 _051_
rlabel metal1 s 1748 18598 1748 18598 4 _052_
rlabel metal2 s 4554 16354 4554 16354 4 _053_
rlabel metal1 s 6532 16762 6532 16762 4 _054_
rlabel metal1 s 6532 14042 6532 14042 4 _055_
rlabel metal1 s 5527 14314 5527 14314 4 _056_
rlabel metal2 s 7038 8738 7038 8738 4 _057_
rlabel metal1 s 7031 11798 7031 11798 4 _058_
rlabel metal2 s 8970 13022 8970 13022 4 _059_
rlabel metal2 s 8970 9758 8970 9758 4 _060_
rlabel metal1 s 7452 15674 7452 15674 4 _061_
rlabel metal2 s 9154 14110 9154 14110 4 _062_
rlabel metal1 s 9292 18190 9292 18190 4 _063_
rlabel metal2 s 9890 15912 9890 15912 4 _064_
rlabel metal1 s 11224 17306 11224 17306 4 _065_
rlabel metal1 s 11677 18734 11677 18734 4 _066_
rlabel metal1 s 10948 14042 10948 14042 4 _067_
rlabel metal1 s 12052 15674 12052 15674 4 _068_
rlabel metal1 s 11047 10710 11047 10710 4 _069_
rlabel metal2 s 11822 13090 11822 13090 4 _070_
rlabel metal2 s 12926 8228 12926 8228 4 _071_
rlabel metal1 s 9706 8058 9706 8058 4 _072_
rlabel metal1 s 13432 11322 13432 11322 4 _073_
rlabel metal1 s 14398 9146 14398 9146 4 _074_
rlabel metal1 s 13715 15470 13715 15470 4 _075_
rlabel metal1 s 14635 13974 14635 13974 4 _076_
rlabel metal1 s 13616 19686 13616 19686 4 _077_
rlabel metal1 s 15371 17238 15371 17238 4 _078_
rlabel metal2 s 17434 19176 17434 19176 4 _079_
rlabel metal1 s 16659 18666 16659 18666 4 _080_
rlabel metal1 s 17388 16218 17388 16218 4 _081_
rlabel metal1 s 17894 17306 17894 17306 4 _082_
rlabel metal2 s 15962 14552 15962 14552 4 _083_
rlabel metal2 s 18538 14212 18538 14212 4 _084_
rlabel metal1 s 15364 11866 15364 11866 4 _085_
rlabel metal2 s 18446 12648 18446 12648 4 _086_
rlabel metal2 s 17710 10472 17710 10472 4 _087_
rlabel metal1 s 16107 9962 16107 9962 4 _088_
rlabel metal2 s 17434 8296 17434 8296 4 _089_
rlabel metal1 s 18407 9622 18407 9622 4 _090_
rlabel metal2 s 15594 6494 15594 6494 4 _091_
rlabel metal1 s 18400 5882 18400 5882 4 _092_
rlabel metal2 s 12926 7208 12926 7208 4 _093_
rlabel metal2 s 15134 5032 15134 5032 4 _094_
rlabel metal2 s 10718 5848 10718 5848 4 _095_
rlabel metal1 s 13340 4794 13340 4794 4 _096_
rlabel metal2 s 15640 14212 15640 14212 4 _097_
rlabel metal2 s 11638 8364 11638 8364 4 _098_
rlabel metal2 s 2852 8398 2852 8398 4 _099_
rlabel metal1 s 2714 5644 2714 5644 4 _100_
rlabel metal1 s 3082 5338 3082 5338 4 _101_
rlabel metal1 s 3634 6358 3634 6358 4 _102_
rlabel metal1 s 9982 6766 9982 6766 4 _103_
rlabel metal1 s 9798 6290 9798 6290 4 _104_
rlabel metal1 s 5382 5814 5382 5814 4 _105_
rlabel metal1 s 8142 5644 8142 5644 4 _106_
rlabel metal1 s 4600 5678 4600 5678 4 _107_
rlabel metal1 s 7176 7174 7176 7174 4 _108_
rlabel metal1 s 6072 7514 6072 7514 4 _109_
rlabel metal1 s 8326 7854 8326 7854 4 _110_
rlabel metal1 s 2438 8534 2438 8534 4 _111_
rlabel metal1 s 2162 8058 2162 8058 4 _112_
rlabel metal1 s 3542 8500 3542 8500 4 _113_
rlabel metal2 s 2346 10608 2346 10608 4 _114_
rlabel metal2 s 3082 11492 3082 11492 4 _115_
rlabel metal2 s 3266 9724 3266 9724 4 _116_
rlabel metal2 s 4554 12852 4554 12852 4 _117_
rlabel metal1 s 5612 11662 5612 11662 4 _118_
rlabel metal1 s 4002 10540 4002 10540 4 _119_
rlabel metal1 s 2392 14450 2392 14450 4 _120_
rlabel metal2 s 2806 14654 2806 14654 4 _121_
rlabel metal2 s 10166 19142 10166 19142 4 _122_
rlabel metal1 s 2599 13906 2599 13906 4 _123_
rlabel metal1 s 3082 18190 3082 18190 4 _124_
rlabel metal1 s 4324 18938 4324 18938 4 _125_
rlabel metal1 s 2898 17204 2898 17204 4 _126_
rlabel metal1 s 5382 18836 5382 18836 4 _127_
rlabel metal1 s 6578 18700 6578 18700 4 _128_
rlabel metal1 s 4554 18394 4554 18394 4 _129_
rlabel metal1 s 4830 17204 4830 17204 4 _130_
rlabel metal1 s 5336 16150 5336 16150 4 _131_
rlabel metal1 s 5697 17170 5697 17170 4 _132_
rlabel metal2 s 12650 11356 12650 11356 4 _133_
rlabel metal1 s 7084 14450 7084 14450 4 _134_
rlabel metal2 s 7498 13668 7498 13668 4 _135_
rlabel metal1 s 6762 15028 6762 15028 4 _136_
rlabel metal2 s 6670 10642 6670 10642 4 _137_
rlabel metal1 s 7682 10166 7682 10166 4 _138_
rlabel metal1 s 6762 11152 6762 11152 4 _139_
rlabel metal2 s 9752 12580 9752 12580 4 _140_
rlabel metal2 s 9338 12818 9338 12818 4 _141_
rlabel metal1 s 8556 11730 8556 11730 4 _142_
rlabel metal1 s 8096 16966 8096 16966 4 _143_
rlabel metal2 s 8326 16388 8326 16388 4 _144_
rlabel metal1 s 8142 15504 8142 15504 4 _145_
rlabel metal1 s 8602 18802 8602 18802 4 _146_
rlabel metal1 s 9660 18734 9660 18734 4 _147_
rlabel metal1 s 8510 18156 8510 18156 4 _148_
rlabel metal1 s 10258 18156 10258 18156 4 _149_
rlabel metal2 s 11086 17612 11086 17612 4 _150_
rlabel metal1 s 9982 19380 9982 19380 4 _151_
rlabel metal1 s 10718 14892 10718 14892 4 _152_
rlabel metal1 s 11638 14042 11638 14042 4 _153_
rlabel metal1 s 16330 14960 16330 14960 4 _154_
rlabel metal1 s 11086 16082 11086 16082 4 _155_
rlabel metal1 s 10580 10234 10580 10234 4 _156_
rlabel metal1 s 11362 10778 11362 10778 4 _157_
rlabel metal1 s 10994 12818 10994 12818 4 _158_
rlabel metal2 s 13386 9282 13386 9282 4 _159_
rlabel metal1 s 13294 8908 13294 8908 4 _160_
rlabel metal1 s 11178 8942 11178 8942 4 _161_
rlabel metal1 s 12466 11254 12466 11254 4 _162_
rlabel metal1 s 12742 11186 12742 11186 4 _163_
rlabel metal1 s 12650 10642 12650 10642 4 _164_
rlabel metal2 s 15870 16796 15870 16796 4 _165_
rlabel metal1 s 13294 14892 13294 14892 4 _166_
rlabel metal1 s 13938 14926 13938 14926 4 _167_
rlabel metal1 s 13570 14450 13570 14450 4 _168_
rlabel metal1 s 13294 18836 13294 18836 4 _169_
rlabel metal1 s 13892 18734 13892 18734 4 _170_
rlabel metal2 s 13386 17850 13386 17850 4 _171_
rlabel metal1 s 17204 18802 17204 18802 4 _172_
rlabel metal1 s 18262 18190 18262 18190 4 _173_
rlabel metal1 s 15364 18258 15364 18258 4 _174_
rlabel metal1 s 17112 17102 17112 17102 4 _175_
rlabel metal1 s 17250 16150 17250 16150 4 _176_
rlabel metal1 s 15916 17170 15916 17170 4 _177_
rlabel metal1 s 17434 13362 17434 13362 4 _178_
rlabel metal1 s 17066 13906 17066 13906 4 _179_
rlabel metal1 s 16744 13294 16744 13294 4 _180_
rlabel metal1 s 16100 12682 16100 12682 4 _181_
rlabel metal2 s 15778 12308 15778 12308 4 _182_
rlabel metal1 s 17066 12614 17066 12614 4 _183_
rlabel metal1 s 16652 10098 16652 10098 4 _184_
rlabel metal1 s 17296 10030 17296 10030 4 _185_
rlabel metal1 s 15226 10676 15226 10676 4 _186_
rlabel metal1 s 16330 8364 16330 8364 4 _187_
rlabel metal2 s 18538 8058 18538 8058 4 _188_
rlabel metal2 s 15870 8500 15870 8500 4 _189_
rlabel metal1 s 16146 5814 16146 5814 4 _190_
rlabel metal1 s 16744 6358 16744 6358 4 _191_
rlabel metal1 s 16790 5746 16790 5746 4 _192_
rlabel metal1 s 15364 7310 15364 7310 4 _193_
rlabel metal1 s 15318 7820 15318 7820 4 _194_
rlabel metal1 s 15410 6766 15410 6766 4 _195_
rlabel metal2 s 11730 5678 11730 5678 4 _196_
rlabel metal1 s 12926 5882 12926 5882 4 _197_
rlabel metal2 s 12650 6154 12650 6154 4 _198_
rlabel metal1 s 14996 8466 14996 8466 4 _199_
rlabel metal1 s 2438 5678 2438 5678 4 _200_
rlabel metal1 s 1794 18836 1794 18836 4 _201_
rlabel metal1 s 6026 13872 6026 13872 4 _202_
rlabel metal1 s 11270 17170 11270 17170 4 _203_
rlabel metal1 s 13938 16048 13938 16048 4 _204_
rlabel metal1 s 18446 13940 18446 13940 4 _205_
rlabel metal2 s 11086 11679 11086 11679 4 clk
rlabel metal1 s 2668 12818 2668 12818 4 clknet_0_clk
rlabel metal2 s 1794 4862 1794 4862 4 clknet_3_0__leaf_clk
rlabel metal1 s 9154 8500 9154 8500 4 clknet_3_1__leaf_clk
rlabel metal1 s 4370 19346 4370 19346 4 clknet_3_2__leaf_clk
rlabel metal1 s 6486 16116 6486 16116 4 clknet_3_3__leaf_clk
rlabel metal2 s 11546 10030 11546 10030 4 clknet_3_4__leaf_clk
rlabel metal1 s 14352 10098 14352 10098 4 clknet_3_5__leaf_clk
rlabel metal1 s 10672 18802 10672 18802 4 clknet_3_6__leaf_clk
rlabel metal1 s 16744 17714 16744 17714 4 clknet_3_7__leaf_clk
rlabel metal1 s 3266 6188 3266 6188 4 csa0.hsum2
rlabel metal1 s 4186 4692 4186 4692 4 csa0.sc
rlabel metal1 s 5244 4658 5244 4658 4 csa0.y
rlabel metal1 s 5290 14450 5290 14450 4 genblk1\[10\].csa.hsum2
rlabel metal2 s 8142 13532 8142 13532 4 genblk1\[10\].csa.sc
rlabel metal2 s 5566 15334 5566 15334 4 genblk1\[10\].csa.sum
rlabel metal2 s 8142 12036 8142 12036 4 genblk1\[10\].csa.y
rlabel metal1 s 6578 11322 6578 11322 4 genblk1\[11\].csa.hsum2
rlabel metal1 s 7728 9554 7728 9554 4 genblk1\[11\].csa.sc
rlabel metal1 s 8142 9418 8142 9418 4 genblk1\[11\].csa.y
rlabel metal2 s 9430 10608 9430 10608 4 genblk1\[12\].csa.hsum2
rlabel metal1 s 10212 12818 10212 12818 4 genblk1\[12\].csa.sc
rlabel metal2 s 10074 13226 10074 13226 4 genblk1\[12\].csa.y
rlabel metal1 s 8687 13702 8687 13702 4 genblk1\[13\].csa.hsum2
rlabel metal2 s 8234 16439 8234 16439 4 genblk1\[13\].csa.sc
rlabel metal1 s 9246 16218 9246 16218 4 genblk1\[13\].csa.y
rlabel metal1 s 10442 16184 10442 16184 4 genblk1\[14\].csa.hsum2
rlabel metal1 s 9522 19346 9522 19346 4 genblk1\[14\].csa.sc
rlabel metal1 s 11270 18292 11270 18292 4 genblk1\[14\].csa.y
rlabel metal1 s 10432 18938 10432 18938 4 genblk1\[15\].csa.hsum2
rlabel metal1 s 12374 17238 12374 17238 4 genblk1\[15\].csa.sc
rlabel metal2 s 12834 16694 12834 16694 4 genblk1\[15\].csa.y
rlabel metal1 s 11362 15980 11362 15980 4 genblk1\[16\].csa.hsum2
rlabel metal1 s 12006 14450 12006 14450 4 genblk1\[16\].csa.sc
rlabel metal1 s 12696 13498 12696 13498 4 genblk1\[16\].csa.y
rlabel metal2 s 11086 13090 11086 13090 4 genblk1\[17\].csa.hsum2
rlabel metal2 s 11086 10914 11086 10914 4 genblk1\[17\].csa.sc
rlabel metal1 s 11592 10030 11592 10030 4 genblk1\[17\].csa.y
rlabel metal1 s 9430 8568 9430 8568 4 genblk1\[18\].csa.hsum2
rlabel metal1 s 13662 8942 13662 8942 4 genblk1\[18\].csa.sc
rlabel metal1 s 13294 9350 13294 9350 4 genblk1\[18\].csa.y
rlabel metal1 s 14168 9486 14168 9486 4 genblk1\[19\].csa.hsum2
rlabel metal1 s 13800 11866 13800 11866 4 genblk1\[19\].csa.sc
rlabel metal1 s 14490 11662 14490 11662 4 genblk1\[19\].csa.y
rlabel metal1 s 4738 5304 4738 5304 4 genblk1\[1\].csa.hsum2
rlabel metal1 s 8602 5675 8602 5675 4 genblk1\[1\].csa.sc
rlabel metal1 s 8924 6222 8924 6222 4 genblk1\[1\].csa.y
rlabel metal1 s 13248 13838 13248 13838 4 genblk1\[20\].csa.hsum2
rlabel metal1 s 14260 15538 14260 15538 4 genblk1\[20\].csa.sc
rlabel metal1 s 15456 15470 15456 15470 4 genblk1\[20\].csa.y
rlabel metal1 s 13938 17272 13938 17272 4 genblk1\[21\].csa.hsum2
rlabel metal1 s 14260 19278 14260 19278 4 genblk1\[21\].csa.sc
rlabel metal1 s 15548 18938 15548 18938 4 genblk1\[21\].csa.y
rlabel metal1 s 15134 18394 15134 18394 4 genblk1\[22\].csa.hsum2
rlabel metal1 s 18400 18802 18400 18802 4 genblk1\[22\].csa.sc
rlabel metal1 s 18722 18292 18722 18292 4 genblk1\[22\].csa.y
rlabel metal1 s 16698 17306 16698 17306 4 genblk1\[23\].csa.hsum2
rlabel metal1 s 18446 16626 18446 16626 4 genblk1\[23\].csa.sc
rlabel metal1 s 18768 16014 18768 16014 4 genblk1\[23\].csa.y
rlabel metal1 s 17250 13498 17250 13498 4 genblk1\[24\].csa.hsum2
rlabel metal1 s 17158 14586 17158 14586 4 genblk1\[24\].csa.sc
rlabel metal1 s 18216 13906 18216 13906 4 genblk1\[24\].csa.y
rlabel metal1 s 17572 12342 17572 12342 4 genblk1\[25\].csa.hsum2
rlabel metal1 s 16146 12274 16146 12274 4 genblk1\[25\].csa.sc
rlabel metal1 s 16008 11730 16008 11730 4 genblk1\[25\].csa.y
rlabel metal1 s 14720 10098 14720 10098 4 genblk1\[26\].csa.hsum2
rlabel metal1 s 18400 10778 18400 10778 4 genblk1\[26\].csa.sc
rlabel metal1 s 18446 10098 18446 10098 4 genblk1\[26\].csa.y
rlabel metal1 s 16192 9146 16192 9146 4 genblk1\[27\].csa.hsum2
rlabel metal1 s 18400 7922 18400 7922 4 genblk1\[27\].csa.sc
rlabel metal1 s 18768 7378 18768 7378 4 genblk1\[27\].csa.y
rlabel metal1 s 17250 5882 17250 5882 4 genblk1\[28\].csa.hsum2
rlabel metal1 s 16606 6154 16606 6154 4 genblk1\[28\].csa.sc
rlabel metal2 s 16330 6018 16330 6018 4 genblk1\[28\].csa.y
rlabel metal1 s 14720 5134 14720 5134 4 genblk1\[29\].csa.hsum2
rlabel metal1 s 13892 7514 13892 7514 4 genblk1\[29\].csa.sc
rlabel metal2 s 14122 6324 14122 6324 4 genblk1\[29\].csa.y
rlabel metal1 s 7544 6358 7544 6358 4 genblk1\[2\].csa.hsum2
rlabel metal1 s 6946 7378 6946 7378 4 genblk1\[2\].csa.sc
rlabel metal1 s 6348 7310 6348 7310 4 genblk1\[2\].csa.y
rlabel metal1 s 12604 5270 12604 5270 4 genblk1\[30\].csa.hsum2
rlabel metal1 s 13386 5780 13386 5780 4 genblk1\[30\].csa.sc
rlabel metal1 s 11178 5338 11178 5338 4 genblk1\[30\].csa.y
rlabel metal1 s 3910 8364 3910 8364 4 genblk1\[3\].csa.hsum2
rlabel metal1 s 2162 8398 2162 8398 4 genblk1\[3\].csa.sc
rlabel metal1 s 1702 9010 1702 9010 4 genblk1\[3\].csa.y
rlabel metal2 s 2898 9826 2898 9826 4 genblk1\[4\].csa.hsum2
rlabel metal1 s 3082 12070 3082 12070 4 genblk1\[4\].csa.sc
rlabel metal2 s 5014 11220 5014 11220 4 genblk1\[4\].csa.y
rlabel metal1 s 4370 10098 4370 10098 4 genblk1\[5\].csa.hsum2
rlabel metal1 s 5336 13294 5336 13294 4 genblk1\[5\].csa.sc
rlabel metal2 s 6210 13158 6210 13158 4 genblk1\[5\].csa.y
rlabel metal2 s 4278 13294 4278 13294 4 genblk1\[6\].csa.hsum2
rlabel metal2 s 3174 15300 3174 15300 4 genblk1\[6\].csa.sc
rlabel metal2 s 3450 15266 3450 15266 4 genblk1\[6\].csa.y
rlabel metal2 s 2898 16796 2898 16796 4 genblk1\[7\].csa.hsum2
rlabel metal1 s 3772 18870 3772 18870 4 genblk1\[7\].csa.sc
rlabel metal1 s 3450 18190 3450 18190 4 genblk1\[7\].csa.y
rlabel metal1 s 2898 18360 2898 18360 4 genblk1\[8\].csa.hsum2
rlabel metal1 s 6440 18802 6440 18802 4 genblk1\[8\].csa.sc
rlabel metal1 s 7406 17850 7406 17850 4 genblk1\[8\].csa.y
rlabel metal1 s 5796 17034 5796 17034 4 genblk1\[9\].csa.hsum2
rlabel metal2 s 5566 16320 5566 16320 4 genblk1\[9\].csa.sc
rlabel metal1 s 15410 2618 15410 2618 4 net1
rlabel metal2 s 11362 16116 11362 16116 4 net10
rlabel metal2 s 11868 16116 11868 16116 4 net11
rlabel metal1 s 12558 11084 12558 11084 4 net12
rlabel metal1 s 2300 19686 2300 19686 4 net13
rlabel metal1 s 13432 14994 13432 14994 4 net14
rlabel metal1 s 13570 18802 13570 18802 4 net15
rlabel metal1 s 14950 19686 14950 19686 4 net16
rlabel metal1 s 15410 17646 15410 17646 4 net17
rlabel metal1 s 16146 15028 16146 15028 4 net18
rlabel metal1 s 15548 12818 15548 12818 4 net19
rlabel metal2 s 2622 6290 2622 6290 4 net2
rlabel metal1 s 15962 10642 15962 10642 4 net20
rlabel metal2 s 17940 13260 17940 13260 4 net21
rlabel metal2 s 17342 19788 17342 19788 4 net22
rlabel metal1 s 15686 7888 15686 7888 4 net23
rlabel metal2 s 4462 16660 4462 16660 4 net24
rlabel metal2 s 18308 16524 18308 16524 4 net25
rlabel metal2 s 18722 16053 18722 16053 4 net26
rlabel metal1 s 3910 8466 3910 8466 4 net27
rlabel metal2 s 2852 16524 2852 16524 4 net28
rlabel metal2 s 4692 12716 4692 12716 4 net29
rlabel metal1 s 7222 15062 7222 15062 4 net3
rlabel metal1 s 2622 14348 2622 14348 4 net30
rlabel metal2 s 3082 19329 3082 19329 4 net31
rlabel metal1 s 5474 18836 5474 18836 4 net32
rlabel metal1 s 6624 19686 6624 19686 4 net33
rlabel metal1 s 1748 16150 1748 16150 4 net34
rlabel metal1 s 1472 5678 1472 5678 4 net35
rlabel metal1 s 9844 7378 9844 7378 4 net36
rlabel metal1 s 7452 9894 7452 9894 4 net37
rlabel metal1 s 7038 10030 7038 10030 4 net38
rlabel metal1 s 9200 5678 9200 5678 4 net39
rlabel metal2 s 7360 16524 7360 16524 4 net4
rlabel metal1 s 5106 5644 5106 5644 4 net40
rlabel metal1 s 8740 16762 8740 16762 4 net41
rlabel metal1 s 8004 16558 8004 16558 4 net42
rlabel metal1 s 13202 5644 13202 5644 4 net43
rlabel metal1 s 12098 6222 12098 6222 4 net44
rlabel metal2 s 4462 10948 4462 10948 4 net45
rlabel metal1 s 2714 11662 2714 11662 4 net46
rlabel metal1 s 14812 19482 14812 19482 4 net47
rlabel metal1 s 10304 18394 10304 18394 4 net48
rlabel metal1 s 8786 18734 8786 18734 4 net49
rlabel metal2 s 9200 13260 9200 13260 4 net5
rlabel metal2 s 7682 12614 7682 12614 4 net50
rlabel metal1 s 6946 14926 6946 14926 4 net51
rlabel metal1 s 14996 19414 14996 19414 4 net52
rlabel metal1 s 7866 12886 7866 12886 4 net53
rlabel metal1 s 16882 11798 16882 11798 4 net54
rlabel metal1 s 17802 12274 17802 12274 4 net55
rlabel metal1 s 11822 13974 11822 13974 4 net56
rlabel metal1 s 11270 14926 11270 14926 4 net57
rlabel metal1 s 7084 9554 7084 9554 4 net58
rlabel metal1 s 13754 12070 13754 12070 4 net59
rlabel metal1 s 8326 16626 8326 16626 4 net6
rlabel metal1 s 14076 8942 14076 8942 4 net60
rlabel metal1 s 12696 9146 12696 9146 4 net61
rlabel metal1 s 6164 11662 6164 11662 4 net62
rlabel metal1 s 4830 11662 4830 11662 4 net63
rlabel metal1 s 3588 5134 3588 5134 4 net64
rlabel metal1 s 14168 7922 14168 7922 4 net65
rlabel metal1 s 11592 10574 11592 10574 4 net66
rlabel metal1 s 14766 7310 14766 7310 4 net67
rlabel metal1 s 4784 18802 4784 18802 4 net68
rlabel metal1 s 17020 6290 17020 6290 4 net69
rlabel metal1 s 9292 18258 9292 18258 4 net7
rlabel metal1 s 16468 6766 16468 6766 4 net70
rlabel metal1 s 12926 17204 12926 17204 4 net71
rlabel metal1 s 6026 16082 6026 16082 4 net72
rlabel metal1 s 7544 18802 7544 18802 4 net73
rlabel metal1 s 5796 18734 5796 18734 4 net74
rlabel metal1 s 3726 14994 3726 14994 4 net75
rlabel metal1 s 9660 13294 9660 13294 4 net76
rlabel metal1 s 1610 7922 1610 7922 4 net77
rlabel metal2 s 2990 8602 2990 8602 4 net78
rlabel metal2 s 18906 10812 18906 10812 4 net79
rlabel metal1 s 10626 19414 10626 19414 4 net8
rlabel metal1 s 18124 13838 18124 13838 4 net80
rlabel metal1 s 15456 15538 15456 15538 4 net81
rlabel metal1 s 7590 7378 7590 7378 4 net82
rlabel metal1 s 18170 16082 18170 16082 4 net83
rlabel metal1 s 11086 10098 11086 10098 4 net84
rlabel metal1 s 19090 18258 19090 18258 4 net85
rlabel metal1 s 19090 7378 19090 7378 4 net86
rlabel metal1 s 11868 10234 11868 10234 4 net87
rlabel metal1 s 14122 6970 14122 6970 4 net88
rlabel metal1 s 10948 15470 10948 15470 4 net9
rlabel metal3 s 1142 5508 1142 5508 4 p
rlabel metal2 s 15226 1027 15226 1027 4 rst
rlabel metal2 s 10350 7650 10350 7650 4 tcmp.z
rlabel metal1 s 1656 19822 1656 19822 4 x[0]
rlabel metal1 s 7268 19822 7268 19822 4 x[10]
rlabel metal1 s 7820 19822 7820 19822 4 x[11]
rlabel metal2 s 8280 19822 8280 19822 4 x[12]
rlabel metal1 s 8970 19822 8970 19822 4 x[13]
rlabel metal1 s 9476 19822 9476 19822 4 x[14]
rlabel metal1 s 9936 19822 9936 19822 4 x[15]
rlabel metal1 s 10488 19822 10488 19822 4 x[16]
rlabel metal2 s 11040 19822 11040 19822 4 x[17]
rlabel metal1 s 11592 19822 11592 19822 4 x[18]
rlabel metal1 s 12144 19822 12144 19822 4 x[19]
rlabel metal1 s 2208 19822 2208 19822 4 x[1]
rlabel metal1 s 12696 19822 12696 19822 4 x[20]
rlabel metal1 s 13938 19856 13938 19856 4 x[21]
rlabel metal1 s 14674 19890 14674 19890 4 x[22]
rlabel metal1 s 14950 19788 14950 19788 4 x[23]
rlabel metal2 s 15180 19822 15180 19822 4 x[24]
rlabel metal1 s 15456 19822 15456 19822 4 x[25]
rlabel metal1 s 16008 19822 16008 19822 4 x[26]
rlabel metal2 s 17526 20094 17526 20094 4 x[27]
rlabel metal1 s 17802 19788 17802 19788 4 x[28]
rlabel metal1 s 18078 19856 18078 19856 4 x[29]
rlabel metal2 s 2714 20818 2714 20818 4 x[2]
rlabel metal1 s 18308 19822 18308 19822 4 x[30]
rlabel metal1 s 18814 19822 18814 19822 4 x[31]
rlabel metal1 s 3220 19822 3220 19822 4 x[3]
rlabel metal1 s 3956 19822 3956 19822 4 x[4]
rlabel metal1 s 4416 19822 4416 19822 4 x[5]
rlabel metal1 s 5060 19822 5060 19822 4 x[6]
rlabel metal1 s 5658 19822 5658 19822 4 x[7]
rlabel metal1 s 6302 19822 6302 19822 4 x[8]
rlabel metal1 s 6854 19856 6854 19856 4 x[9]
rlabel metal3 s 820 16660 820 16660 4 y
flabel metal5 s 1056 18384 19276 18704 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 13896 19276 14216 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 9408 19276 9728 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4920 19276 5240 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 17462 2128 17782 20176 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12931 2128 13251 20176 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8400 2128 8720 20176 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3869 2128 4189 20176 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 17724 19276 18044 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 13236 19276 13556 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8748 19276 9068 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4260 19276 4580 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 16802 2128 17122 20176 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12271 2128 12591 20176 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7740 2128 8060 20176 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3209 2128 3529 20176 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 19570 11160 20370 11280 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 p
port 4 nsew
flabel metal2 s 15198 0 15254 800 0 FreeSans 280 90 0 0 rst
port 5 nsew
flabel metal2 s 1582 21714 1638 22514 0 FreeSans 280 90 0 0 x[0]
port 6 nsew
flabel metal2 s 7102 21714 7158 22514 0 FreeSans 280 90 0 0 x[10]
port 7 nsew
flabel metal2 s 7654 21714 7710 22514 0 FreeSans 280 90 0 0 x[11]
port 8 nsew
flabel metal2 s 8206 21714 8262 22514 0 FreeSans 280 90 0 0 x[12]
port 9 nsew
flabel metal2 s 8758 21714 8814 22514 0 FreeSans 280 90 0 0 x[13]
port 10 nsew
flabel metal2 s 9310 21714 9366 22514 0 FreeSans 280 90 0 0 x[14]
port 11 nsew
flabel metal2 s 9862 21714 9918 22514 0 FreeSans 280 90 0 0 x[15]
port 12 nsew
flabel metal2 s 10414 21714 10470 22514 0 FreeSans 280 90 0 0 x[16]
port 13 nsew
flabel metal2 s 10966 21714 11022 22514 0 FreeSans 280 90 0 0 x[17]
port 14 nsew
flabel metal2 s 11518 21714 11574 22514 0 FreeSans 280 90 0 0 x[18]
port 15 nsew
flabel metal2 s 12070 21714 12126 22514 0 FreeSans 280 90 0 0 x[19]
port 16 nsew
flabel metal2 s 2134 21714 2190 22514 0 FreeSans 280 90 0 0 x[1]
port 17 nsew
flabel metal2 s 12622 21714 12678 22514 0 FreeSans 280 90 0 0 x[20]
port 18 nsew
flabel metal2 s 13174 21714 13230 22514 0 FreeSans 280 90 0 0 x[21]
port 19 nsew
flabel metal2 s 13726 21714 13782 22514 0 FreeSans 280 90 0 0 x[22]
port 20 nsew
flabel metal2 s 14278 21714 14334 22514 0 FreeSans 280 90 0 0 x[23]
port 21 nsew
flabel metal2 s 14830 21714 14886 22514 0 FreeSans 280 90 0 0 x[24]
port 22 nsew
flabel metal2 s 15382 21714 15438 22514 0 FreeSans 280 90 0 0 x[25]
port 23 nsew
flabel metal2 s 15934 21714 15990 22514 0 FreeSans 280 90 0 0 x[26]
port 24 nsew
flabel metal2 s 16486 21714 16542 22514 0 FreeSans 280 90 0 0 x[27]
port 25 nsew
flabel metal2 s 17038 21714 17094 22514 0 FreeSans 280 90 0 0 x[28]
port 26 nsew
flabel metal2 s 17590 21714 17646 22514 0 FreeSans 280 90 0 0 x[29]
port 27 nsew
flabel metal2 s 2686 21714 2742 22514 0 FreeSans 280 90 0 0 x[2]
port 28 nsew
flabel metal2 s 18142 21714 18198 22514 0 FreeSans 280 90 0 0 x[30]
port 29 nsew
flabel metal2 s 18694 21714 18750 22514 0 FreeSans 280 90 0 0 x[31]
port 30 nsew
flabel metal2 s 3238 21714 3294 22514 0 FreeSans 280 90 0 0 x[3]
port 31 nsew
flabel metal2 s 3790 21714 3846 22514 0 FreeSans 280 90 0 0 x[4]
port 32 nsew
flabel metal2 s 4342 21714 4398 22514 0 FreeSans 280 90 0 0 x[5]
port 33 nsew
flabel metal2 s 4894 21714 4950 22514 0 FreeSans 280 90 0 0 x[6]
port 34 nsew
flabel metal2 s 5446 21714 5502 22514 0 FreeSans 280 90 0 0 x[7]
port 35 nsew
flabel metal2 s 5998 21714 6054 22514 0 FreeSans 280 90 0 0 x[8]
port 36 nsew
flabel metal2 s 6550 21714 6606 22514 0 FreeSans 280 90 0 0 x[9]
port 37 nsew
flabel metal3 s 0 16600 800 16720 0 FreeSans 600 0 0 0 y
port 38 nsew
<< properties >>
string FIXED_BBOX 0 0 20370 22514
<< end >>
